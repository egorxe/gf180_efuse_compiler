VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array
  CLASS BLOCK ;
  FOREIGN efuse_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 193.820 BY 60.305 ;
  PIN COL_PROG[0]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 178.440 59.415 178.780 60.305 ;
    END
  END COL_PROG[0]
  PIN COL_PROG[1]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 183.080 59.415 183.420 60.305 ;
    END
  END COL_PROG[1]
  PIN COL_PROG[2]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 187.720 59.415 188.060 60.305 ;
    END
  END COL_PROG[2]
  PIN COL_PROG[3]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 192.360 59.415 192.700 60.305 ;
    END
  END COL_PROG[3]
  PIN DO[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.720 1.770 17.100 2.150 ;
        RECT 16.745 0.000 17.075 1.770 ;
    END
  END DO[0]
  PIN LINE[0]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 18.305 2.770 18.685 3.150 ;
        RECT 18.330 0.000 18.660 2.770 ;
    END
  END LINE[0]
  PIN DO[1]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.910 1.770 35.290 2.150 ;
        RECT 34.935 0.000 35.265 1.770 ;
    END
  END DO[1]
  PIN LINE[1]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 36.495 2.770 36.875 3.150 ;
        RECT 36.520 0.000 36.850 2.770 ;
    END
  END LINE[1]
  PIN DO[2]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.220 1.770 54.600 2.150 ;
        RECT 54.245 0.000 54.575 1.770 ;
    END
  END DO[2]
  PIN DO[3]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.050 1.770 69.430 2.150 ;
        RECT 69.075 0.000 69.405 1.770 ;
    END
  END DO[3]
  PIN LINE[2]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 70.635 2.770 71.015 3.150 ;
        RECT 70.660 0.000 70.990 2.770 ;
    END
  END LINE[2]
  PIN LINE[3]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 79.595 2.770 79.975 3.150 ;
        RECT 79.620 0.000 79.950 2.770 ;
    END
  END LINE[3]
  PIN LINE[4]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 101.995 2.770 102.375 3.150 ;
        RECT 102.020 0.000 102.350 2.770 ;
    END
  END LINE[4]
  PIN LINE[5]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 122.155 2.770 122.535 3.150 ;
        RECT 122.180 0.000 122.510 2.770 ;
    END
  END LINE[5]
  PIN LINE[6]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 144.555 2.770 144.935 3.150 ;
        RECT 144.580 0.000 144.910 2.770 ;
    END
  END LINE[6]
  PIN LINE[7]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 166.955 2.770 167.335 3.150 ;
        RECT 166.980 0.000 167.310 2.770 ;
    END
  END LINE[7]
  PIN SENSE
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER Metal3 ;
        RECT 4.170 3.775 4.550 3.800 ;
        RECT 22.360 3.775 22.740 3.800 ;
        RECT 41.670 3.775 42.050 3.800 ;
        RECT 56.500 3.775 56.880 3.800 ;
        RECT 4.170 3.445 56.880 3.775 ;
        RECT 4.170 3.420 4.550 3.445 ;
        RECT 22.360 3.420 22.740 3.445 ;
        RECT 41.670 3.420 42.050 3.445 ;
        RECT 56.500 3.420 56.880 3.445 ;
    END
  END SENSE
  PIN nPRESET
    ANTENNAGATEAREA 3.800000 ;
    PORT
      LAYER Metal3 ;
        RECT 4.580 3.115 4.960 3.140 ;
        RECT 22.770 3.115 23.150 3.140 ;
        RECT 42.080 3.115 42.460 3.140 ;
        RECT 56.910 3.115 57.290 3.140 ;
        RECT 4.580 2.785 57.290 3.115 ;
        RECT 4.580 2.760 4.960 2.785 ;
        RECT 22.770 2.760 23.150 2.785 ;
        RECT 42.080 2.760 42.460 2.785 ;
        RECT 56.910 2.760 57.290 2.785 ;
    END
  END nPRESET
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 57.805 193.820 60.305 ;
        RECT 0.000 49.035 1.910 57.805 ;
        RECT 10.290 49.035 12.200 57.805 ;
        RECT 20.575 49.035 23.905 57.805 ;
        RECT 32.285 49.035 34.195 57.805 ;
        RECT 42.570 49.035 45.900 57.805 ;
        RECT 54.280 49.035 56.190 57.805 ;
        RECT 64.565 49.035 67.895 57.805 ;
        RECT 76.275 49.035 78.185 57.805 ;
        RECT 86.560 49.035 89.890 57.805 ;
        RECT 98.270 49.035 100.180 57.805 ;
        RECT 108.555 49.035 111.885 57.805 ;
        RECT 120.265 49.035 122.175 57.805 ;
        RECT 130.550 49.035 133.880 57.805 ;
        RECT 142.260 49.035 144.170 57.805 ;
        RECT 152.545 49.035 155.875 57.805 ;
        RECT 164.255 49.035 166.165 57.805 ;
        RECT 173.540 49.035 176.450 57.805 ;
        RECT 173.540 6.470 176.040 49.035 ;
        RECT 0.000 3.970 176.040 6.470 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 177.175 55.495 179.290 55.805 ;
        RECT 181.815 55.495 183.930 55.805 ;
        RECT 186.455 55.495 188.570 55.805 ;
        RECT 191.095 55.495 193.210 55.805 ;
        RECT 177.150 55.115 179.315 55.495 ;
        RECT 181.790 55.115 183.955 55.495 ;
        RECT 186.430 55.115 188.595 55.495 ;
        RECT 191.070 55.115 193.235 55.495 ;
        RECT 177.175 54.835 179.290 55.115 ;
        RECT 181.815 54.835 183.930 55.115 ;
        RECT 186.455 54.835 188.570 55.115 ;
        RECT 191.095 54.835 193.210 55.115 ;
        RECT 177.150 54.455 179.315 54.835 ;
        RECT 181.790 54.455 183.955 54.835 ;
        RECT 186.430 54.455 188.595 54.835 ;
        RECT 191.070 54.455 193.235 54.835 ;
        RECT 177.175 54.175 179.290 54.455 ;
        RECT 181.815 54.175 183.930 54.455 ;
        RECT 186.455 54.175 188.570 54.455 ;
        RECT 191.095 54.175 193.210 54.455 ;
        RECT 177.150 53.795 179.315 54.175 ;
        RECT 181.790 53.795 183.955 54.175 ;
        RECT 186.430 53.795 188.595 54.175 ;
        RECT 191.070 53.795 193.235 54.175 ;
        RECT 177.175 53.515 179.290 53.795 ;
        RECT 181.815 53.515 183.930 53.795 ;
        RECT 186.455 53.515 188.570 53.795 ;
        RECT 191.095 53.515 193.210 53.795 ;
        RECT 177.150 53.135 179.315 53.515 ;
        RECT 181.790 53.135 183.955 53.515 ;
        RECT 186.430 53.135 188.595 53.515 ;
        RECT 191.070 53.135 193.235 53.515 ;
        RECT 177.175 52.855 179.290 53.135 ;
        RECT 181.815 52.855 183.930 53.135 ;
        RECT 186.455 52.855 188.570 53.135 ;
        RECT 191.095 52.855 193.210 53.135 ;
        RECT 177.150 52.475 179.315 52.855 ;
        RECT 181.790 52.475 183.955 52.855 ;
        RECT 186.430 52.475 188.595 52.855 ;
        RECT 191.070 52.475 193.235 52.855 ;
        RECT 177.175 52.195 179.290 52.475 ;
        RECT 181.815 52.195 183.930 52.475 ;
        RECT 186.455 52.195 188.570 52.475 ;
        RECT 191.095 52.195 193.210 52.475 ;
        RECT 177.150 51.815 179.315 52.195 ;
        RECT 181.790 51.815 183.955 52.195 ;
        RECT 186.430 51.815 188.595 52.195 ;
        RECT 191.070 51.815 193.235 52.195 ;
        RECT 177.175 51.535 179.290 51.815 ;
        RECT 181.815 51.535 183.930 51.815 ;
        RECT 186.455 51.535 188.570 51.815 ;
        RECT 191.095 51.535 193.210 51.815 ;
        RECT 177.150 51.155 179.315 51.535 ;
        RECT 181.790 51.155 183.955 51.535 ;
        RECT 186.430 51.155 188.595 51.535 ;
        RECT 191.070 51.155 193.235 51.535 ;
        RECT 177.175 50.875 179.290 51.155 ;
        RECT 181.815 50.875 183.930 51.155 ;
        RECT 186.455 50.875 188.570 51.155 ;
        RECT 191.095 50.875 193.210 51.155 ;
        RECT 177.150 50.495 179.315 50.875 ;
        RECT 181.790 50.495 183.955 50.875 ;
        RECT 186.430 50.495 188.595 50.875 ;
        RECT 191.070 50.495 193.235 50.875 ;
        RECT 177.175 18.495 179.290 50.495 ;
        RECT 181.815 18.495 183.930 50.495 ;
        RECT 186.455 18.495 188.570 50.495 ;
        RECT 191.095 18.495 193.210 50.495 ;
        RECT 177.150 18.115 179.315 18.495 ;
        RECT 181.790 18.115 183.955 18.495 ;
        RECT 186.430 18.115 188.595 18.495 ;
        RECT 191.070 18.115 193.235 18.495 ;
        RECT 177.175 17.835 179.290 18.115 ;
        RECT 181.815 17.835 183.930 18.115 ;
        RECT 186.455 17.835 188.570 18.115 ;
        RECT 191.095 17.835 193.210 18.115 ;
        RECT 177.150 17.455 179.315 17.835 ;
        RECT 181.790 17.455 183.955 17.835 ;
        RECT 186.430 17.455 188.595 17.835 ;
        RECT 191.070 17.455 193.235 17.835 ;
        RECT 177.175 17.175 179.290 17.455 ;
        RECT 181.815 17.175 183.930 17.455 ;
        RECT 186.455 17.175 188.570 17.455 ;
        RECT 191.095 17.175 193.210 17.455 ;
        RECT 177.150 16.795 179.315 17.175 ;
        RECT 181.790 16.795 183.955 17.175 ;
        RECT 186.430 16.795 188.595 17.175 ;
        RECT 191.070 16.795 193.235 17.175 ;
        RECT 177.175 16.515 179.290 16.795 ;
        RECT 181.815 16.515 183.930 16.795 ;
        RECT 186.455 16.515 188.570 16.795 ;
        RECT 191.095 16.515 193.210 16.795 ;
        RECT 177.150 16.135 179.315 16.515 ;
        RECT 181.790 16.135 183.955 16.515 ;
        RECT 186.430 16.135 188.595 16.515 ;
        RECT 191.070 16.135 193.235 16.515 ;
        RECT 177.175 15.855 179.290 16.135 ;
        RECT 181.815 15.855 183.930 16.135 ;
        RECT 186.455 15.855 188.570 16.135 ;
        RECT 191.095 15.855 193.210 16.135 ;
        RECT 177.150 15.475 179.315 15.855 ;
        RECT 181.790 15.475 183.955 15.855 ;
        RECT 186.430 15.475 188.595 15.855 ;
        RECT 191.070 15.475 193.235 15.855 ;
        RECT 177.175 15.195 179.290 15.475 ;
        RECT 181.815 15.195 183.930 15.475 ;
        RECT 186.455 15.195 188.570 15.475 ;
        RECT 191.095 15.195 193.210 15.475 ;
        RECT 177.150 14.815 179.315 15.195 ;
        RECT 181.790 14.815 183.955 15.195 ;
        RECT 186.430 14.815 188.595 15.195 ;
        RECT 191.070 14.815 193.235 15.195 ;
        RECT 177.175 14.535 179.290 14.815 ;
        RECT 181.815 14.535 183.930 14.815 ;
        RECT 186.455 14.535 188.570 14.815 ;
        RECT 191.095 14.535 193.210 14.815 ;
        RECT 177.150 14.155 179.315 14.535 ;
        RECT 181.790 14.155 183.955 14.535 ;
        RECT 186.430 14.155 188.595 14.535 ;
        RECT 191.070 14.155 193.235 14.535 ;
        RECT 177.175 13.875 179.290 14.155 ;
        RECT 181.815 13.875 183.930 14.155 ;
        RECT 186.455 13.875 188.570 14.155 ;
        RECT 191.095 13.875 193.210 14.155 ;
        RECT 177.150 13.495 179.315 13.875 ;
        RECT 181.790 13.495 183.955 13.875 ;
        RECT 186.430 13.495 188.595 13.875 ;
        RECT 191.070 13.495 193.235 13.875 ;
        RECT 177.175 13.215 179.290 13.495 ;
        RECT 181.815 13.215 183.930 13.495 ;
        RECT 186.455 13.215 188.570 13.495 ;
        RECT 191.095 13.215 193.210 13.495 ;
        RECT 177.150 12.835 179.315 13.215 ;
        RECT 181.790 12.835 183.955 13.215 ;
        RECT 186.430 12.835 188.595 13.215 ;
        RECT 191.070 12.835 193.235 13.215 ;
        RECT 177.175 12.555 179.290 12.835 ;
        RECT 181.815 12.555 183.930 12.835 ;
        RECT 186.455 12.555 188.570 12.835 ;
        RECT 191.095 12.555 193.210 12.835 ;
        RECT 177.150 12.175 179.315 12.555 ;
        RECT 181.790 12.175 183.955 12.555 ;
        RECT 186.430 12.175 188.595 12.555 ;
        RECT 191.070 12.175 193.235 12.555 ;
        RECT 177.175 11.895 179.290 12.175 ;
        RECT 181.815 11.895 183.930 12.175 ;
        RECT 186.455 11.895 188.570 12.175 ;
        RECT 191.095 11.895 193.210 12.175 ;
        RECT 177.150 11.515 179.315 11.895 ;
        RECT 181.790 11.515 183.955 11.895 ;
        RECT 186.430 11.515 188.595 11.895 ;
        RECT 191.070 11.515 193.235 11.895 ;
        RECT 177.175 11.235 179.290 11.515 ;
        RECT 181.815 11.235 183.930 11.515 ;
        RECT 186.455 11.235 188.570 11.515 ;
        RECT 191.095 11.235 193.210 11.515 ;
        RECT 177.150 10.855 179.315 11.235 ;
        RECT 181.790 10.855 183.955 11.235 ;
        RECT 186.430 10.855 188.595 11.235 ;
        RECT 191.070 10.855 193.235 11.235 ;
        RECT 177.175 10.575 179.290 10.855 ;
        RECT 181.815 10.575 183.930 10.855 ;
        RECT 186.455 10.575 188.570 10.855 ;
        RECT 191.095 10.575 193.210 10.855 ;
        RECT 177.150 10.195 179.315 10.575 ;
        RECT 181.790 10.195 183.955 10.575 ;
        RECT 186.430 10.195 188.595 10.575 ;
        RECT 191.070 10.195 193.235 10.575 ;
        RECT 177.175 9.915 179.290 10.195 ;
        RECT 181.815 9.915 183.930 10.195 ;
        RECT 186.455 9.915 188.570 10.195 ;
        RECT 191.095 9.915 193.210 10.195 ;
        RECT 177.150 9.535 179.315 9.915 ;
        RECT 181.790 9.535 183.955 9.915 ;
        RECT 186.430 9.535 188.595 9.915 ;
        RECT 191.070 9.535 193.235 9.915 ;
        RECT 177.175 9.255 179.290 9.535 ;
        RECT 181.815 9.255 183.930 9.535 ;
        RECT 186.455 9.255 188.570 9.535 ;
        RECT 191.095 9.255 193.210 9.535 ;
        RECT 177.150 8.875 179.315 9.255 ;
        RECT 181.790 8.875 183.955 9.255 ;
        RECT 186.430 8.875 188.595 9.255 ;
        RECT 191.070 8.875 193.235 9.255 ;
        RECT 177.175 2.500 179.290 8.875 ;
        RECT 181.815 2.500 183.930 8.875 ;
        RECT 186.455 2.500 188.570 8.875 ;
        RECT 191.095 2.500 193.210 8.875 ;
        RECT 0.000 0.000 193.820 2.500 ;
    END
  END VDD
  OBS
      LAYER Metal1 ;
        RECT 1.975 59.605 2.675 60.305 ;
        RECT 0.735 9.370 1.905 59.380 ;
        RECT 1.525 9.360 1.905 9.370 ;
        RECT 2.755 56.865 6.970 59.380 ;
        RECT 2.755 9.360 3.125 56.865 ;
        RECT 5.220 54.845 6.970 56.865 ;
        RECT 5.690 49.385 6.500 53.395 ;
        RECT 5.250 46.485 6.950 49.385 ;
        RECT 5.250 19.685 6.950 22.585 ;
        RECT 5.700 15.660 6.510 19.685 ;
        RECT 5.230 12.190 6.980 14.210 ;
        RECT 9.075 12.190 9.445 59.695 ;
        RECT 5.230 9.675 9.445 12.190 ;
        RECT 10.295 59.685 10.675 59.695 ;
        RECT 11.815 59.685 12.195 59.695 ;
        RECT 10.295 9.675 12.195 59.685 ;
        RECT 13.045 12.190 13.415 59.695 ;
        RECT 19.810 59.605 20.510 60.305 ;
        RECT 23.970 59.605 24.670 60.305 ;
        RECT 15.515 56.865 19.730 59.380 ;
        RECT 15.515 54.845 17.265 56.865 ;
        RECT 15.985 49.385 16.795 53.395 ;
        RECT 15.550 43.785 17.250 49.385 ;
        RECT 15.550 19.685 17.250 25.285 ;
        RECT 15.980 15.660 16.790 19.685 ;
        RECT 15.510 12.190 17.260 14.210 ;
        RECT 13.045 9.675 17.260 12.190 ;
        RECT 9.525 8.750 10.225 9.450 ;
        RECT 12.265 8.750 12.965 9.450 ;
        RECT 19.360 9.360 19.730 56.865 ;
        RECT 20.580 9.370 21.750 59.380 ;
        RECT 22.730 9.370 23.900 59.380 ;
        RECT 20.580 9.360 20.960 9.370 ;
        RECT 23.520 9.360 23.900 9.370 ;
        RECT 24.750 56.865 28.965 59.380 ;
        RECT 24.750 9.360 25.120 56.865 ;
        RECT 27.215 54.845 28.965 56.865 ;
        RECT 27.685 49.385 28.495 53.395 ;
        RECT 27.245 46.485 28.945 49.385 ;
        RECT 27.245 19.685 28.945 22.585 ;
        RECT 27.695 15.660 28.505 19.685 ;
        RECT 27.225 12.190 28.975 14.210 ;
        RECT 31.070 12.190 31.440 59.695 ;
        RECT 27.225 9.675 31.440 12.190 ;
        RECT 32.290 59.685 32.670 59.695 ;
        RECT 33.810 59.685 34.190 59.695 ;
        RECT 32.290 9.675 34.190 59.685 ;
        RECT 35.040 12.190 35.410 59.695 ;
        RECT 41.805 59.605 42.505 60.305 ;
        RECT 45.965 59.605 46.665 60.305 ;
        RECT 37.510 56.865 41.725 59.380 ;
        RECT 37.510 54.845 39.260 56.865 ;
        RECT 37.980 49.385 38.790 53.395 ;
        RECT 37.545 43.785 39.245 49.385 ;
        RECT 37.545 19.685 39.245 25.285 ;
        RECT 37.975 15.660 38.785 19.685 ;
        RECT 37.505 12.190 39.255 14.210 ;
        RECT 35.040 9.675 39.255 12.190 ;
        RECT 31.520 8.750 32.220 9.450 ;
        RECT 34.260 8.750 34.960 9.450 ;
        RECT 41.355 9.360 41.725 56.865 ;
        RECT 42.575 9.370 43.745 59.380 ;
        RECT 44.725 9.370 45.895 59.380 ;
        RECT 42.575 9.360 42.955 9.370 ;
        RECT 45.515 9.360 45.895 9.370 ;
        RECT 46.745 56.865 50.960 59.380 ;
        RECT 46.745 9.360 47.115 56.865 ;
        RECT 49.210 54.845 50.960 56.865 ;
        RECT 49.680 49.385 50.490 53.395 ;
        RECT 49.240 46.485 50.940 49.385 ;
        RECT 49.240 19.685 50.940 22.585 ;
        RECT 49.690 15.660 50.500 19.685 ;
        RECT 49.220 12.190 50.970 14.210 ;
        RECT 53.065 12.190 53.435 59.695 ;
        RECT 49.220 9.675 53.435 12.190 ;
        RECT 54.285 59.685 54.665 59.695 ;
        RECT 55.805 59.685 56.185 59.695 ;
        RECT 54.285 9.675 56.185 59.685 ;
        RECT 57.035 12.190 57.405 59.695 ;
        RECT 63.800 59.605 64.500 60.305 ;
        RECT 67.960 59.605 68.660 60.305 ;
        RECT 59.505 56.865 63.720 59.380 ;
        RECT 59.505 54.845 61.255 56.865 ;
        RECT 59.975 49.385 60.785 53.395 ;
        RECT 59.540 43.785 61.240 49.385 ;
        RECT 59.540 19.685 61.240 25.285 ;
        RECT 59.970 15.660 60.780 19.685 ;
        RECT 59.500 12.190 61.250 14.210 ;
        RECT 57.035 9.675 61.250 12.190 ;
        RECT 53.515 8.750 54.215 9.450 ;
        RECT 56.255 8.750 56.955 9.450 ;
        RECT 63.350 9.360 63.720 56.865 ;
        RECT 64.570 9.370 65.740 59.380 ;
        RECT 66.720 9.370 67.890 59.380 ;
        RECT 64.570 9.360 64.950 9.370 ;
        RECT 67.510 9.360 67.890 9.370 ;
        RECT 68.740 56.865 72.955 59.380 ;
        RECT 68.740 9.360 69.110 56.865 ;
        RECT 71.205 54.845 72.955 56.865 ;
        RECT 71.675 49.385 72.485 53.395 ;
        RECT 71.235 46.485 72.935 49.385 ;
        RECT 71.235 19.685 72.935 22.585 ;
        RECT 71.685 15.660 72.495 19.685 ;
        RECT 71.215 12.190 72.965 14.210 ;
        RECT 75.060 12.190 75.430 59.695 ;
        RECT 71.215 9.675 75.430 12.190 ;
        RECT 76.280 59.685 76.660 59.695 ;
        RECT 77.800 59.685 78.180 59.695 ;
        RECT 76.280 9.675 78.180 59.685 ;
        RECT 79.030 12.190 79.400 59.695 ;
        RECT 85.795 59.605 86.495 60.305 ;
        RECT 89.955 59.605 90.655 60.305 ;
        RECT 81.500 56.865 85.715 59.380 ;
        RECT 81.500 54.845 83.250 56.865 ;
        RECT 81.970 49.385 82.780 53.395 ;
        RECT 81.535 43.785 83.235 49.385 ;
        RECT 81.535 19.685 83.235 25.285 ;
        RECT 81.965 15.660 82.775 19.685 ;
        RECT 81.495 12.190 83.245 14.210 ;
        RECT 79.030 9.675 83.245 12.190 ;
        RECT 75.510 8.750 76.210 9.450 ;
        RECT 78.250 8.750 78.950 9.450 ;
        RECT 85.345 9.360 85.715 56.865 ;
        RECT 86.565 9.370 87.735 59.380 ;
        RECT 88.715 9.370 89.885 59.380 ;
        RECT 86.565 9.360 86.945 9.370 ;
        RECT 89.505 9.360 89.885 9.370 ;
        RECT 90.735 56.865 94.950 59.380 ;
        RECT 90.735 9.360 91.105 56.865 ;
        RECT 93.200 54.845 94.950 56.865 ;
        RECT 93.670 49.385 94.480 53.395 ;
        RECT 93.230 46.485 94.930 49.385 ;
        RECT 93.230 19.685 94.930 22.585 ;
        RECT 93.680 15.660 94.490 19.685 ;
        RECT 93.210 12.190 94.960 14.210 ;
        RECT 97.055 12.190 97.425 59.695 ;
        RECT 93.210 9.675 97.425 12.190 ;
        RECT 98.275 59.685 98.655 59.695 ;
        RECT 99.795 59.685 100.175 59.695 ;
        RECT 98.275 9.675 100.175 59.685 ;
        RECT 101.025 12.190 101.395 59.695 ;
        RECT 107.790 59.605 108.490 60.305 ;
        RECT 111.950 59.605 112.650 60.305 ;
        RECT 103.495 56.865 107.710 59.380 ;
        RECT 103.495 54.845 105.245 56.865 ;
        RECT 103.965 49.385 104.775 53.395 ;
        RECT 103.530 43.785 105.230 49.385 ;
        RECT 103.530 19.685 105.230 25.285 ;
        RECT 103.960 15.660 104.770 19.685 ;
        RECT 103.490 12.190 105.240 14.210 ;
        RECT 101.025 9.675 105.240 12.190 ;
        RECT 97.505 8.750 98.205 9.450 ;
        RECT 100.245 8.750 100.945 9.450 ;
        RECT 107.340 9.360 107.710 56.865 ;
        RECT 108.560 9.370 109.730 59.380 ;
        RECT 110.710 9.370 111.880 59.380 ;
        RECT 108.560 9.360 108.940 9.370 ;
        RECT 111.500 9.360 111.880 9.370 ;
        RECT 112.730 56.865 116.945 59.380 ;
        RECT 112.730 9.360 113.100 56.865 ;
        RECT 115.195 54.845 116.945 56.865 ;
        RECT 115.665 49.385 116.475 53.395 ;
        RECT 115.225 46.485 116.925 49.385 ;
        RECT 115.225 19.685 116.925 22.585 ;
        RECT 115.675 15.660 116.485 19.685 ;
        RECT 115.205 12.190 116.955 14.210 ;
        RECT 119.050 12.190 119.420 59.695 ;
        RECT 115.205 9.675 119.420 12.190 ;
        RECT 120.270 59.685 120.650 59.695 ;
        RECT 121.790 59.685 122.170 59.695 ;
        RECT 120.270 9.675 122.170 59.685 ;
        RECT 123.020 12.190 123.390 59.695 ;
        RECT 129.785 59.605 130.485 60.305 ;
        RECT 133.945 59.605 134.645 60.305 ;
        RECT 125.490 56.865 129.705 59.380 ;
        RECT 125.490 54.845 127.240 56.865 ;
        RECT 125.960 49.385 126.770 53.395 ;
        RECT 125.525 43.785 127.225 49.385 ;
        RECT 125.525 19.685 127.225 25.285 ;
        RECT 125.955 15.660 126.765 19.685 ;
        RECT 125.485 12.190 127.235 14.210 ;
        RECT 123.020 9.675 127.235 12.190 ;
        RECT 119.500 8.750 120.200 9.450 ;
        RECT 122.240 8.750 122.940 9.450 ;
        RECT 129.335 9.360 129.705 56.865 ;
        RECT 130.555 9.370 131.725 59.380 ;
        RECT 132.705 9.370 133.875 59.380 ;
        RECT 130.555 9.360 130.935 9.370 ;
        RECT 133.495 9.360 133.875 9.370 ;
        RECT 134.725 56.865 138.940 59.380 ;
        RECT 134.725 9.360 135.095 56.865 ;
        RECT 137.190 54.845 138.940 56.865 ;
        RECT 137.660 49.385 138.470 53.395 ;
        RECT 137.220 46.485 138.920 49.385 ;
        RECT 137.220 19.685 138.920 22.585 ;
        RECT 137.670 15.660 138.480 19.685 ;
        RECT 137.200 12.190 138.950 14.210 ;
        RECT 141.045 12.190 141.415 59.695 ;
        RECT 137.200 9.675 141.415 12.190 ;
        RECT 142.265 59.685 142.645 59.695 ;
        RECT 143.785 59.685 144.165 59.695 ;
        RECT 142.265 9.675 144.165 59.685 ;
        RECT 145.015 12.190 145.385 59.695 ;
        RECT 151.780 59.605 152.480 60.305 ;
        RECT 155.940 59.605 156.640 60.305 ;
        RECT 147.485 56.865 151.700 59.380 ;
        RECT 147.485 54.845 149.235 56.865 ;
        RECT 147.955 49.385 148.765 53.395 ;
        RECT 147.520 43.785 149.220 49.385 ;
        RECT 147.520 19.685 149.220 25.285 ;
        RECT 147.950 15.660 148.760 19.685 ;
        RECT 147.480 12.190 149.230 14.210 ;
        RECT 145.015 9.675 149.230 12.190 ;
        RECT 141.495 8.750 142.195 9.450 ;
        RECT 144.235 8.750 144.935 9.450 ;
        RECT 151.330 9.360 151.700 56.865 ;
        RECT 152.550 9.370 153.720 59.380 ;
        RECT 154.700 9.370 155.870 59.380 ;
        RECT 152.550 9.360 152.930 9.370 ;
        RECT 155.490 9.360 155.870 9.370 ;
        RECT 156.720 56.865 160.935 59.380 ;
        RECT 156.720 9.360 157.090 56.865 ;
        RECT 159.185 54.845 160.935 56.865 ;
        RECT 159.655 49.385 160.465 53.395 ;
        RECT 159.215 46.485 160.915 49.385 ;
        RECT 159.215 19.685 160.915 22.585 ;
        RECT 159.665 15.660 160.475 19.685 ;
        RECT 159.195 12.190 160.945 14.210 ;
        RECT 163.040 12.190 163.410 59.695 ;
        RECT 159.195 9.675 163.410 12.190 ;
        RECT 164.260 59.685 164.640 59.695 ;
        RECT 165.780 59.685 166.160 59.695 ;
        RECT 164.260 9.675 166.160 59.685 ;
        RECT 167.010 12.190 167.380 59.695 ;
        RECT 173.775 59.605 174.475 60.305 ;
        RECT 169.480 56.865 173.695 59.380 ;
        RECT 169.480 54.845 171.230 56.865 ;
        RECT 169.950 49.385 170.760 53.395 ;
        RECT 169.515 43.785 171.215 49.385 ;
        RECT 169.515 19.685 171.215 25.285 ;
        RECT 169.945 15.660 170.755 19.685 ;
        RECT 169.475 12.190 171.225 14.210 ;
        RECT 167.010 9.675 171.225 12.190 ;
        RECT 163.490 8.750 164.190 9.450 ;
        RECT 166.230 8.750 166.930 9.450 ;
        RECT 173.325 9.360 173.695 56.865 ;
        RECT 174.545 9.370 175.715 59.380 ;
        RECT 174.545 9.360 174.925 9.370 ;
        RECT 177.120 9.185 177.560 59.185 ;
        RECT 177.150 8.875 177.530 9.185 ;
        RECT 177.910 9.175 178.290 59.195 ;
        RECT 178.940 55.495 179.310 59.195 ;
        RECT 178.935 55.115 179.315 55.495 ;
        RECT 178.940 54.835 179.310 55.115 ;
        RECT 178.935 54.455 179.315 54.835 ;
        RECT 178.940 54.175 179.310 54.455 ;
        RECT 178.935 53.795 179.315 54.175 ;
        RECT 178.940 53.515 179.310 53.795 ;
        RECT 178.935 53.135 179.315 53.515 ;
        RECT 178.940 52.855 179.310 53.135 ;
        RECT 178.935 52.475 179.315 52.855 ;
        RECT 178.940 52.195 179.310 52.475 ;
        RECT 178.935 51.815 179.315 52.195 ;
        RECT 178.940 51.535 179.310 51.815 ;
        RECT 178.935 51.155 179.315 51.535 ;
        RECT 178.940 50.875 179.310 51.155 ;
        RECT 178.935 50.495 179.315 50.875 ;
        RECT 178.940 18.495 179.310 50.495 ;
        RECT 178.935 18.115 179.315 18.495 ;
        RECT 178.940 17.835 179.310 18.115 ;
        RECT 178.935 17.455 179.315 17.835 ;
        RECT 178.940 17.175 179.310 17.455 ;
        RECT 178.935 16.795 179.315 17.175 ;
        RECT 178.940 16.515 179.310 16.795 ;
        RECT 178.935 16.135 179.315 16.515 ;
        RECT 178.940 15.855 179.310 16.135 ;
        RECT 178.935 15.475 179.315 15.855 ;
        RECT 178.940 15.195 179.310 15.475 ;
        RECT 178.935 14.815 179.315 15.195 ;
        RECT 178.940 14.535 179.310 14.815 ;
        RECT 178.935 14.155 179.315 14.535 ;
        RECT 178.940 13.875 179.310 14.155 ;
        RECT 178.935 13.495 179.315 13.875 ;
        RECT 178.940 13.215 179.310 13.495 ;
        RECT 178.935 12.835 179.315 13.215 ;
        RECT 178.940 12.555 179.310 12.835 ;
        RECT 178.935 12.175 179.315 12.555 ;
        RECT 178.940 11.895 179.310 12.175 ;
        RECT 178.935 11.515 179.315 11.895 ;
        RECT 178.940 11.235 179.310 11.515 ;
        RECT 178.935 10.855 179.315 11.235 ;
        RECT 178.940 10.575 179.310 10.855 ;
        RECT 178.935 10.195 179.315 10.575 ;
        RECT 178.940 9.915 179.310 10.195 ;
        RECT 178.935 9.535 179.315 9.915 ;
        RECT 178.940 9.255 179.310 9.535 ;
        RECT 178.935 8.875 179.315 9.255 ;
        RECT 181.760 9.185 182.200 59.185 ;
        RECT 181.790 8.875 182.170 9.185 ;
        RECT 182.550 9.175 182.930 59.195 ;
        RECT 183.580 55.495 183.950 59.195 ;
        RECT 183.575 55.115 183.955 55.495 ;
        RECT 183.580 54.835 183.950 55.115 ;
        RECT 183.575 54.455 183.955 54.835 ;
        RECT 183.580 54.175 183.950 54.455 ;
        RECT 183.575 53.795 183.955 54.175 ;
        RECT 183.580 53.515 183.950 53.795 ;
        RECT 183.575 53.135 183.955 53.515 ;
        RECT 183.580 52.855 183.950 53.135 ;
        RECT 183.575 52.475 183.955 52.855 ;
        RECT 183.580 52.195 183.950 52.475 ;
        RECT 183.575 51.815 183.955 52.195 ;
        RECT 183.580 51.535 183.950 51.815 ;
        RECT 183.575 51.155 183.955 51.535 ;
        RECT 183.580 50.875 183.950 51.155 ;
        RECT 183.575 50.495 183.955 50.875 ;
        RECT 183.580 18.495 183.950 50.495 ;
        RECT 183.575 18.115 183.955 18.495 ;
        RECT 183.580 17.835 183.950 18.115 ;
        RECT 183.575 17.455 183.955 17.835 ;
        RECT 183.580 17.175 183.950 17.455 ;
        RECT 183.575 16.795 183.955 17.175 ;
        RECT 183.580 16.515 183.950 16.795 ;
        RECT 183.575 16.135 183.955 16.515 ;
        RECT 183.580 15.855 183.950 16.135 ;
        RECT 183.575 15.475 183.955 15.855 ;
        RECT 183.580 15.195 183.950 15.475 ;
        RECT 183.575 14.815 183.955 15.195 ;
        RECT 183.580 14.535 183.950 14.815 ;
        RECT 183.575 14.155 183.955 14.535 ;
        RECT 183.580 13.875 183.950 14.155 ;
        RECT 183.575 13.495 183.955 13.875 ;
        RECT 183.580 13.215 183.950 13.495 ;
        RECT 183.575 12.835 183.955 13.215 ;
        RECT 183.580 12.555 183.950 12.835 ;
        RECT 183.575 12.175 183.955 12.555 ;
        RECT 183.580 11.895 183.950 12.175 ;
        RECT 183.575 11.515 183.955 11.895 ;
        RECT 183.580 11.235 183.950 11.515 ;
        RECT 183.575 10.855 183.955 11.235 ;
        RECT 183.580 10.575 183.950 10.855 ;
        RECT 183.575 10.195 183.955 10.575 ;
        RECT 183.580 9.915 183.950 10.195 ;
        RECT 183.575 9.535 183.955 9.915 ;
        RECT 183.580 9.255 183.950 9.535 ;
        RECT 183.575 8.875 183.955 9.255 ;
        RECT 186.400 9.185 186.840 59.185 ;
        RECT 186.430 8.875 186.810 9.185 ;
        RECT 187.190 9.175 187.570 59.195 ;
        RECT 188.220 55.495 188.590 59.195 ;
        RECT 188.215 55.115 188.595 55.495 ;
        RECT 188.220 54.835 188.590 55.115 ;
        RECT 188.215 54.455 188.595 54.835 ;
        RECT 188.220 54.175 188.590 54.455 ;
        RECT 188.215 53.795 188.595 54.175 ;
        RECT 188.220 53.515 188.590 53.795 ;
        RECT 188.215 53.135 188.595 53.515 ;
        RECT 188.220 52.855 188.590 53.135 ;
        RECT 188.215 52.475 188.595 52.855 ;
        RECT 188.220 52.195 188.590 52.475 ;
        RECT 188.215 51.815 188.595 52.195 ;
        RECT 188.220 51.535 188.590 51.815 ;
        RECT 188.215 51.155 188.595 51.535 ;
        RECT 188.220 50.875 188.590 51.155 ;
        RECT 188.215 50.495 188.595 50.875 ;
        RECT 188.220 18.495 188.590 50.495 ;
        RECT 188.215 18.115 188.595 18.495 ;
        RECT 188.220 17.835 188.590 18.115 ;
        RECT 188.215 17.455 188.595 17.835 ;
        RECT 188.220 17.175 188.590 17.455 ;
        RECT 188.215 16.795 188.595 17.175 ;
        RECT 188.220 16.515 188.590 16.795 ;
        RECT 188.215 16.135 188.595 16.515 ;
        RECT 188.220 15.855 188.590 16.135 ;
        RECT 188.215 15.475 188.595 15.855 ;
        RECT 188.220 15.195 188.590 15.475 ;
        RECT 188.215 14.815 188.595 15.195 ;
        RECT 188.220 14.535 188.590 14.815 ;
        RECT 188.215 14.155 188.595 14.535 ;
        RECT 188.220 13.875 188.590 14.155 ;
        RECT 188.215 13.495 188.595 13.875 ;
        RECT 188.220 13.215 188.590 13.495 ;
        RECT 188.215 12.835 188.595 13.215 ;
        RECT 188.220 12.555 188.590 12.835 ;
        RECT 188.215 12.175 188.595 12.555 ;
        RECT 188.220 11.895 188.590 12.175 ;
        RECT 188.215 11.515 188.595 11.895 ;
        RECT 188.220 11.235 188.590 11.515 ;
        RECT 188.215 10.855 188.595 11.235 ;
        RECT 188.220 10.575 188.590 10.855 ;
        RECT 188.215 10.195 188.595 10.575 ;
        RECT 188.220 9.915 188.590 10.195 ;
        RECT 188.215 9.535 188.595 9.915 ;
        RECT 188.220 9.255 188.590 9.535 ;
        RECT 188.215 8.875 188.595 9.255 ;
        RECT 191.040 9.185 191.480 59.185 ;
        RECT 191.070 8.875 191.450 9.185 ;
        RECT 191.830 9.175 192.210 59.195 ;
        RECT 192.860 55.495 193.230 59.195 ;
        RECT 192.855 55.115 193.235 55.495 ;
        RECT 192.860 54.835 193.230 55.115 ;
        RECT 192.855 54.455 193.235 54.835 ;
        RECT 192.860 54.175 193.230 54.455 ;
        RECT 192.855 53.795 193.235 54.175 ;
        RECT 192.860 53.515 193.230 53.795 ;
        RECT 192.855 53.135 193.235 53.515 ;
        RECT 192.860 52.855 193.230 53.135 ;
        RECT 192.855 52.475 193.235 52.855 ;
        RECT 192.860 52.195 193.230 52.475 ;
        RECT 192.855 51.815 193.235 52.195 ;
        RECT 192.860 51.535 193.230 51.815 ;
        RECT 192.855 51.155 193.235 51.535 ;
        RECT 192.860 50.875 193.230 51.155 ;
        RECT 192.855 50.495 193.235 50.875 ;
        RECT 192.860 18.495 193.230 50.495 ;
        RECT 192.855 18.115 193.235 18.495 ;
        RECT 192.860 17.835 193.230 18.115 ;
        RECT 192.855 17.455 193.235 17.835 ;
        RECT 192.860 17.175 193.230 17.455 ;
        RECT 192.855 16.795 193.235 17.175 ;
        RECT 192.860 16.515 193.230 16.795 ;
        RECT 192.855 16.135 193.235 16.515 ;
        RECT 192.860 15.855 193.230 16.135 ;
        RECT 192.855 15.475 193.235 15.855 ;
        RECT 192.860 15.195 193.230 15.475 ;
        RECT 192.855 14.815 193.235 15.195 ;
        RECT 192.860 14.535 193.230 14.815 ;
        RECT 192.855 14.155 193.235 14.535 ;
        RECT 192.860 13.875 193.230 14.155 ;
        RECT 192.855 13.495 193.235 13.875 ;
        RECT 192.860 13.215 193.230 13.495 ;
        RECT 192.855 12.835 193.235 13.215 ;
        RECT 192.860 12.555 193.230 12.835 ;
        RECT 192.855 12.175 193.235 12.555 ;
        RECT 192.860 11.895 193.230 12.175 ;
        RECT 192.855 11.515 193.235 11.895 ;
        RECT 192.860 11.235 193.230 11.515 ;
        RECT 192.855 10.855 193.235 11.235 ;
        RECT 192.860 10.575 193.230 10.855 ;
        RECT 192.855 10.195 193.235 10.575 ;
        RECT 192.860 9.915 193.230 10.195 ;
        RECT 192.855 9.535 193.235 9.915 ;
        RECT 192.860 9.255 193.230 9.535 ;
        RECT 192.855 8.875 193.235 9.255 ;
        RECT 0.500 4.580 2.740 5.180 ;
        RECT 0.870 3.690 1.210 4.580 ;
        RECT 2.010 3.695 2.350 4.580 ;
        RECT 3.490 4.030 3.860 4.550 ;
        RECT 4.610 4.030 4.990 8.470 ;
        RECT 5.340 4.580 20.930 5.180 ;
        RECT 5.340 4.040 5.780 4.580 ;
        RECT 4.170 3.740 4.550 3.800 ;
        RECT 3.455 3.420 4.550 3.740 ;
        RECT 6.615 3.720 6.845 4.580 ;
        RECT 3.455 3.410 4.540 3.420 ;
        RECT 0.870 1.260 1.210 2.960 ;
        RECT 2.010 1.260 2.350 2.950 ;
        RECT 4.270 2.820 5.270 3.150 ;
        RECT 4.580 2.760 4.960 2.820 ;
        RECT 7.080 2.680 7.405 3.680 ;
        RECT 7.635 3.330 7.965 4.350 ;
        RECT 8.855 3.720 9.085 4.580 ;
        RECT 9.320 3.330 9.645 3.680 ;
        RECT 7.635 3.065 9.645 3.330 ;
        RECT 0.500 0.660 2.740 1.260 ;
        RECT 3.820 0.610 4.190 2.530 ;
        RECT 4.840 1.260 5.220 2.530 ;
        RECT 5.570 1.260 6.010 2.520 ;
        RECT 6.715 1.260 6.945 2.350 ;
        RECT 7.635 1.490 7.965 3.065 ;
        RECT 9.320 2.680 9.645 3.065 ;
        RECT 8.955 1.260 9.185 2.350 ;
        RECT 9.875 1.490 10.205 4.350 ;
        RECT 11.095 3.930 11.325 4.580 ;
        RECT 12.245 3.660 12.475 4.350 ;
        RECT 13.365 3.930 13.595 4.580 ;
        RECT 12.245 3.405 13.530 3.660 ;
        RECT 11.480 2.760 13.000 3.175 ;
        RECT 13.230 2.520 13.530 3.405 ;
        RECT 11.095 1.260 11.325 2.240 ;
        RECT 12.070 2.200 13.530 2.520 ;
        RECT 14.455 2.300 14.685 4.080 ;
        RECT 14.915 3.250 15.430 4.230 ;
        RECT 15.795 4.015 16.025 4.580 ;
        RECT 16.540 3.280 17.165 4.305 ;
        RECT 14.915 2.690 15.800 3.250 ;
        RECT 16.180 2.300 16.465 3.050 ;
        RECT 12.070 1.490 12.520 2.200 ;
        RECT 14.455 2.065 16.465 2.300 ;
        RECT 13.365 1.260 13.595 1.950 ;
        RECT 14.455 1.490 14.840 2.065 ;
        RECT 15.740 1.260 16.080 1.750 ;
        RECT 16.695 1.500 17.165 3.280 ;
        RECT 17.815 2.300 18.045 4.080 ;
        RECT 18.275 3.250 18.790 4.230 ;
        RECT 19.155 4.015 19.385 4.580 ;
        RECT 19.900 3.280 20.525 4.305 ;
        RECT 21.680 4.030 22.050 4.550 ;
        RECT 22.800 4.030 23.180 8.470 ;
        RECT 23.530 4.580 40.240 5.180 ;
        RECT 23.530 4.040 23.970 4.580 ;
        RECT 22.360 3.740 22.740 3.800 ;
        RECT 21.645 3.420 22.740 3.740 ;
        RECT 24.805 3.720 25.035 4.580 ;
        RECT 21.645 3.410 22.730 3.420 ;
        RECT 18.275 2.690 19.160 3.250 ;
        RECT 19.540 2.300 19.825 3.050 ;
        RECT 17.815 2.065 19.825 2.300 ;
        RECT 17.815 1.490 18.200 2.065 ;
        RECT 19.100 1.260 19.440 1.750 ;
        RECT 20.055 1.500 20.525 3.280 ;
        RECT 22.460 2.820 23.460 3.150 ;
        RECT 22.770 2.760 23.150 2.820 ;
        RECT 25.270 2.680 25.595 3.680 ;
        RECT 25.825 3.330 26.155 4.350 ;
        RECT 27.045 3.720 27.275 4.580 ;
        RECT 27.510 3.330 27.835 3.680 ;
        RECT 25.825 3.065 27.835 3.330 ;
        RECT 4.840 0.660 20.930 1.260 ;
        RECT 4.840 0.610 5.220 0.660 ;
        RECT 5.570 0.620 6.010 0.660 ;
        RECT 22.010 0.610 22.380 2.530 ;
        RECT 23.030 1.260 23.410 2.530 ;
        RECT 23.760 1.260 24.200 2.520 ;
        RECT 24.905 1.260 25.135 2.350 ;
        RECT 25.825 1.490 26.155 3.065 ;
        RECT 27.510 2.680 27.835 3.065 ;
        RECT 27.145 1.260 27.375 2.350 ;
        RECT 28.065 1.490 28.395 4.350 ;
        RECT 29.285 3.930 29.515 4.580 ;
        RECT 30.435 3.660 30.665 4.350 ;
        RECT 31.555 3.930 31.785 4.580 ;
        RECT 30.435 3.405 31.720 3.660 ;
        RECT 29.670 2.760 31.190 3.175 ;
        RECT 31.420 2.520 31.720 3.405 ;
        RECT 29.285 1.260 29.515 2.240 ;
        RECT 30.260 2.200 31.720 2.520 ;
        RECT 32.645 2.300 32.875 4.080 ;
        RECT 33.105 3.250 33.620 4.230 ;
        RECT 33.985 4.015 34.215 4.580 ;
        RECT 34.730 3.280 35.355 4.305 ;
        RECT 33.105 2.690 33.990 3.250 ;
        RECT 34.370 2.300 34.655 3.050 ;
        RECT 30.260 1.490 30.710 2.200 ;
        RECT 32.645 2.065 34.655 2.300 ;
        RECT 31.555 1.260 31.785 1.950 ;
        RECT 32.645 1.490 33.030 2.065 ;
        RECT 33.930 1.260 34.270 1.750 ;
        RECT 34.885 1.500 35.355 3.280 ;
        RECT 36.005 2.300 36.235 4.080 ;
        RECT 36.465 3.250 36.980 4.230 ;
        RECT 37.345 4.015 37.575 4.580 ;
        RECT 38.090 3.280 38.715 4.305 ;
        RECT 39.510 3.695 39.850 4.580 ;
        RECT 40.990 4.030 41.360 4.550 ;
        RECT 42.110 4.030 42.490 8.470 ;
        RECT 42.840 4.580 55.070 5.180 ;
        RECT 42.840 4.040 43.280 4.580 ;
        RECT 41.670 3.740 42.050 3.800 ;
        RECT 40.955 3.420 42.050 3.740 ;
        RECT 44.115 3.720 44.345 4.580 ;
        RECT 40.955 3.410 42.040 3.420 ;
        RECT 36.465 2.690 37.350 3.250 ;
        RECT 37.730 2.300 38.015 3.050 ;
        RECT 36.005 2.065 38.015 2.300 ;
        RECT 36.005 1.490 36.390 2.065 ;
        RECT 37.290 1.260 37.630 1.750 ;
        RECT 38.245 1.500 38.715 3.280 ;
        RECT 39.510 1.260 39.850 2.950 ;
        RECT 41.770 2.820 42.770 3.150 ;
        RECT 42.080 2.760 42.460 2.820 ;
        RECT 44.580 2.680 44.905 3.680 ;
        RECT 45.135 3.330 45.465 4.350 ;
        RECT 46.355 3.720 46.585 4.580 ;
        RECT 46.820 3.330 47.145 3.680 ;
        RECT 45.135 3.065 47.145 3.330 ;
        RECT 23.030 0.660 40.240 1.260 ;
        RECT 23.030 0.610 23.410 0.660 ;
        RECT 23.760 0.620 24.200 0.660 ;
        RECT 41.320 0.610 41.690 2.530 ;
        RECT 42.340 1.260 42.720 2.530 ;
        RECT 43.070 1.260 43.510 2.520 ;
        RECT 44.215 1.260 44.445 2.350 ;
        RECT 45.135 1.490 45.465 3.065 ;
        RECT 46.820 2.680 47.145 3.065 ;
        RECT 46.455 1.260 46.685 2.350 ;
        RECT 47.375 1.490 47.705 4.350 ;
        RECT 48.595 3.930 48.825 4.580 ;
        RECT 49.745 3.660 49.975 4.350 ;
        RECT 50.865 3.930 51.095 4.580 ;
        RECT 49.745 3.405 51.030 3.660 ;
        RECT 48.980 2.760 50.500 3.175 ;
        RECT 50.730 2.520 51.030 3.405 ;
        RECT 48.595 1.260 48.825 2.240 ;
        RECT 49.570 2.200 51.030 2.520 ;
        RECT 51.955 2.300 52.185 4.080 ;
        RECT 52.415 3.250 52.930 4.230 ;
        RECT 53.295 4.015 53.525 4.580 ;
        RECT 54.040 3.280 54.665 4.305 ;
        RECT 55.820 4.030 56.190 4.550 ;
        RECT 56.940 4.030 57.320 8.470 ;
        RECT 57.670 4.580 175.180 5.180 ;
        RECT 57.670 4.040 58.110 4.580 ;
        RECT 56.500 3.740 56.880 3.800 ;
        RECT 55.785 3.420 56.880 3.740 ;
        RECT 58.945 3.720 59.175 4.580 ;
        RECT 55.785 3.410 56.870 3.420 ;
        RECT 52.415 2.690 53.300 3.250 ;
        RECT 53.680 2.300 53.965 3.050 ;
        RECT 49.570 1.490 50.020 2.200 ;
        RECT 51.955 2.065 53.965 2.300 ;
        RECT 50.865 1.260 51.095 1.950 ;
        RECT 51.955 1.490 52.340 2.065 ;
        RECT 53.240 1.260 53.580 1.750 ;
        RECT 54.195 1.500 54.665 3.280 ;
        RECT 56.600 2.820 57.600 3.150 ;
        RECT 56.910 2.760 57.290 2.820 ;
        RECT 59.410 2.680 59.735 3.680 ;
        RECT 59.965 3.330 60.295 4.350 ;
        RECT 61.185 3.720 61.415 4.580 ;
        RECT 61.650 3.330 61.975 3.680 ;
        RECT 59.965 3.065 61.975 3.330 ;
        RECT 42.340 0.660 55.070 1.260 ;
        RECT 42.340 0.610 42.720 0.660 ;
        RECT 43.070 0.620 43.510 0.660 ;
        RECT 56.150 0.610 56.520 2.530 ;
        RECT 57.170 1.260 57.550 2.530 ;
        RECT 57.900 1.260 58.340 2.520 ;
        RECT 59.045 1.260 59.275 2.350 ;
        RECT 59.965 1.490 60.295 3.065 ;
        RECT 61.650 2.680 61.975 3.065 ;
        RECT 61.285 1.260 61.515 2.350 ;
        RECT 62.205 1.490 62.535 4.350 ;
        RECT 63.425 3.930 63.655 4.580 ;
        RECT 64.575 3.660 64.805 4.350 ;
        RECT 65.695 3.930 65.925 4.580 ;
        RECT 64.575 3.405 65.860 3.660 ;
        RECT 63.810 2.760 65.330 3.175 ;
        RECT 65.560 2.520 65.860 3.405 ;
        RECT 63.425 1.260 63.655 2.240 ;
        RECT 64.400 2.200 65.860 2.520 ;
        RECT 66.785 2.300 67.015 4.080 ;
        RECT 67.245 3.250 67.760 4.230 ;
        RECT 68.125 4.015 68.355 4.580 ;
        RECT 68.870 3.280 69.495 4.305 ;
        RECT 67.245 2.690 68.130 3.250 ;
        RECT 68.510 2.300 68.795 3.050 ;
        RECT 64.400 1.490 64.850 2.200 ;
        RECT 66.785 2.065 68.795 2.300 ;
        RECT 65.695 1.260 65.925 1.950 ;
        RECT 66.785 1.490 67.170 2.065 ;
        RECT 68.070 1.260 68.410 1.750 ;
        RECT 69.025 1.500 69.495 3.280 ;
        RECT 70.145 2.300 70.375 4.080 ;
        RECT 70.605 3.250 71.120 4.230 ;
        RECT 71.485 4.015 71.715 4.580 ;
        RECT 72.230 3.280 72.855 4.305 ;
        RECT 73.650 3.695 73.990 4.580 ;
        RECT 74.625 3.785 74.855 4.580 ;
        RECT 70.605 2.690 71.490 3.250 ;
        RECT 71.870 2.300 72.155 3.050 ;
        RECT 70.145 2.065 72.155 2.300 ;
        RECT 70.145 1.490 70.530 2.065 ;
        RECT 71.430 1.260 71.770 1.750 ;
        RECT 72.385 1.500 72.855 3.280 ;
        RECT 74.625 3.325 75.900 3.555 ;
        RECT 73.650 1.260 73.990 2.950 ;
        RECT 74.625 1.490 74.855 3.325 ;
        RECT 76.145 2.920 76.375 4.350 ;
        RECT 76.865 3.785 77.095 4.580 ;
        RECT 75.110 2.690 76.375 2.920 ;
        RECT 76.865 3.325 78.140 3.555 ;
        RECT 76.145 1.260 76.375 2.390 ;
        RECT 76.865 1.490 77.095 3.325 ;
        RECT 78.385 2.920 78.615 4.350 ;
        RECT 77.350 2.690 78.615 2.920 ;
        RECT 78.385 1.260 78.615 2.390 ;
        RECT 79.105 2.300 79.335 4.080 ;
        RECT 79.565 3.250 80.080 4.230 ;
        RECT 80.445 4.015 80.675 4.580 ;
        RECT 81.190 3.280 81.815 4.305 ;
        RECT 82.465 3.785 82.695 4.580 ;
        RECT 79.565 2.690 80.450 3.250 ;
        RECT 80.830 2.300 81.115 3.050 ;
        RECT 79.105 2.065 81.115 2.300 ;
        RECT 79.105 1.490 79.490 2.065 ;
        RECT 80.390 1.260 80.730 1.750 ;
        RECT 81.345 1.500 81.815 3.280 ;
        RECT 82.465 3.325 83.740 3.555 ;
        RECT 82.465 1.490 82.695 3.325 ;
        RECT 83.985 2.920 84.215 4.350 ;
        RECT 84.705 3.785 84.935 4.580 ;
        RECT 82.950 2.690 84.215 2.920 ;
        RECT 84.705 3.325 85.980 3.555 ;
        RECT 83.985 1.260 84.215 2.390 ;
        RECT 84.705 1.490 84.935 3.325 ;
        RECT 86.225 2.920 86.455 4.350 ;
        RECT 86.945 3.785 87.175 4.580 ;
        RECT 85.190 2.690 86.455 2.920 ;
        RECT 86.945 3.325 88.220 3.555 ;
        RECT 86.225 1.260 86.455 2.390 ;
        RECT 86.945 1.490 87.175 3.325 ;
        RECT 88.465 2.920 88.695 4.350 ;
        RECT 89.185 3.785 89.415 4.580 ;
        RECT 87.430 2.690 88.695 2.920 ;
        RECT 89.185 3.325 90.460 3.555 ;
        RECT 88.465 1.260 88.695 2.390 ;
        RECT 89.185 1.490 89.415 3.325 ;
        RECT 90.705 2.920 90.935 4.350 ;
        RECT 91.425 3.785 91.655 4.580 ;
        RECT 89.670 2.690 90.935 2.920 ;
        RECT 91.425 3.325 92.700 3.555 ;
        RECT 90.705 1.260 90.935 2.390 ;
        RECT 91.425 1.490 91.655 3.325 ;
        RECT 92.945 2.920 93.175 4.350 ;
        RECT 93.810 3.695 94.150 4.580 ;
        RECT 94.785 3.785 95.015 4.580 ;
        RECT 94.785 3.325 96.060 3.555 ;
        RECT 91.910 2.690 93.175 2.920 ;
        RECT 92.945 1.260 93.175 2.390 ;
        RECT 93.810 1.260 94.150 2.950 ;
        RECT 94.785 1.490 95.015 3.325 ;
        RECT 96.305 2.920 96.535 4.350 ;
        RECT 97.025 3.785 97.255 4.580 ;
        RECT 95.270 2.690 96.535 2.920 ;
        RECT 97.025 3.325 98.300 3.555 ;
        RECT 96.305 1.260 96.535 2.390 ;
        RECT 97.025 1.490 97.255 3.325 ;
        RECT 98.545 2.920 98.775 4.350 ;
        RECT 99.265 3.785 99.495 4.580 ;
        RECT 97.510 2.690 98.775 2.920 ;
        RECT 99.265 3.325 100.540 3.555 ;
        RECT 98.545 1.260 98.775 2.390 ;
        RECT 99.265 1.490 99.495 3.325 ;
        RECT 100.785 2.920 101.015 4.350 ;
        RECT 99.750 2.690 101.015 2.920 ;
        RECT 100.785 1.260 101.015 2.390 ;
        RECT 101.505 2.300 101.735 4.080 ;
        RECT 101.965 3.250 102.480 4.230 ;
        RECT 102.845 4.015 103.075 4.580 ;
        RECT 103.590 3.280 104.215 4.305 ;
        RECT 104.865 3.785 105.095 4.580 ;
        RECT 101.965 2.690 102.850 3.250 ;
        RECT 103.230 2.300 103.515 3.050 ;
        RECT 101.505 2.065 103.515 2.300 ;
        RECT 101.505 1.490 101.890 2.065 ;
        RECT 102.790 1.260 103.130 1.750 ;
        RECT 103.745 1.500 104.215 3.280 ;
        RECT 104.865 3.325 106.140 3.555 ;
        RECT 104.865 1.490 105.095 3.325 ;
        RECT 106.385 2.920 106.615 4.350 ;
        RECT 107.105 3.785 107.335 4.580 ;
        RECT 105.350 2.690 106.615 2.920 ;
        RECT 107.105 3.325 108.380 3.555 ;
        RECT 106.385 1.260 106.615 2.390 ;
        RECT 107.105 1.490 107.335 3.325 ;
        RECT 108.625 2.920 108.855 4.350 ;
        RECT 109.345 3.785 109.575 4.580 ;
        RECT 107.590 2.690 108.855 2.920 ;
        RECT 109.345 3.325 110.620 3.555 ;
        RECT 108.625 1.260 108.855 2.390 ;
        RECT 109.345 1.490 109.575 3.325 ;
        RECT 110.865 2.920 111.095 4.350 ;
        RECT 111.585 3.785 111.815 4.580 ;
        RECT 109.830 2.690 111.095 2.920 ;
        RECT 111.585 3.325 112.860 3.555 ;
        RECT 110.865 1.260 111.095 2.390 ;
        RECT 111.585 1.490 111.815 3.325 ;
        RECT 113.105 2.920 113.335 4.350 ;
        RECT 113.970 3.695 114.310 4.580 ;
        RECT 114.945 3.785 115.175 4.580 ;
        RECT 114.945 3.325 116.220 3.555 ;
        RECT 112.070 2.690 113.335 2.920 ;
        RECT 113.105 1.260 113.335 2.390 ;
        RECT 113.970 1.260 114.310 2.950 ;
        RECT 114.945 1.490 115.175 3.325 ;
        RECT 116.465 2.920 116.695 4.350 ;
        RECT 117.185 3.785 117.415 4.580 ;
        RECT 115.430 2.690 116.695 2.920 ;
        RECT 117.185 3.325 118.460 3.555 ;
        RECT 116.465 1.260 116.695 2.390 ;
        RECT 117.185 1.490 117.415 3.325 ;
        RECT 118.705 2.920 118.935 4.350 ;
        RECT 119.425 3.785 119.655 4.580 ;
        RECT 117.670 2.690 118.935 2.920 ;
        RECT 119.425 3.325 120.700 3.555 ;
        RECT 118.705 1.260 118.935 2.390 ;
        RECT 119.425 1.490 119.655 3.325 ;
        RECT 120.945 2.920 121.175 4.350 ;
        RECT 119.910 2.690 121.175 2.920 ;
        RECT 120.945 1.260 121.175 2.390 ;
        RECT 121.665 2.300 121.895 4.080 ;
        RECT 122.125 3.250 122.640 4.230 ;
        RECT 123.005 4.015 123.235 4.580 ;
        RECT 123.750 3.280 124.375 4.305 ;
        RECT 125.025 3.785 125.255 4.580 ;
        RECT 122.125 2.690 123.010 3.250 ;
        RECT 123.390 2.300 123.675 3.050 ;
        RECT 121.665 2.065 123.675 2.300 ;
        RECT 121.665 1.490 122.050 2.065 ;
        RECT 122.950 1.260 123.290 1.750 ;
        RECT 123.905 1.500 124.375 3.280 ;
        RECT 125.025 3.325 126.300 3.555 ;
        RECT 125.025 1.490 125.255 3.325 ;
        RECT 126.545 2.920 126.775 4.350 ;
        RECT 127.265 3.785 127.495 4.580 ;
        RECT 125.510 2.690 126.775 2.920 ;
        RECT 127.265 3.325 128.540 3.555 ;
        RECT 126.545 1.260 126.775 2.390 ;
        RECT 127.265 1.490 127.495 3.325 ;
        RECT 128.785 2.920 129.015 4.350 ;
        RECT 129.505 3.785 129.735 4.580 ;
        RECT 127.750 2.690 129.015 2.920 ;
        RECT 129.505 3.325 130.780 3.555 ;
        RECT 128.785 1.260 129.015 2.390 ;
        RECT 129.505 1.490 129.735 3.325 ;
        RECT 131.025 2.920 131.255 4.350 ;
        RECT 131.745 3.785 131.975 4.580 ;
        RECT 129.990 2.690 131.255 2.920 ;
        RECT 131.745 3.325 133.020 3.555 ;
        RECT 131.025 1.260 131.255 2.390 ;
        RECT 131.745 1.490 131.975 3.325 ;
        RECT 133.265 2.920 133.495 4.350 ;
        RECT 134.130 3.695 134.470 4.580 ;
        RECT 135.105 3.785 135.335 4.580 ;
        RECT 135.105 3.325 136.380 3.555 ;
        RECT 132.230 2.690 133.495 2.920 ;
        RECT 133.265 1.260 133.495 2.390 ;
        RECT 134.130 1.260 134.470 2.950 ;
        RECT 135.105 1.490 135.335 3.325 ;
        RECT 136.625 2.920 136.855 4.350 ;
        RECT 137.345 3.785 137.575 4.580 ;
        RECT 135.590 2.690 136.855 2.920 ;
        RECT 137.345 3.325 138.620 3.555 ;
        RECT 136.625 1.260 136.855 2.390 ;
        RECT 137.345 1.490 137.575 3.325 ;
        RECT 138.865 2.920 139.095 4.350 ;
        RECT 139.585 3.785 139.815 4.580 ;
        RECT 137.830 2.690 139.095 2.920 ;
        RECT 139.585 3.325 140.860 3.555 ;
        RECT 138.865 1.260 139.095 2.390 ;
        RECT 139.585 1.490 139.815 3.325 ;
        RECT 141.105 2.920 141.335 4.350 ;
        RECT 141.825 3.785 142.055 4.580 ;
        RECT 140.070 2.690 141.335 2.920 ;
        RECT 141.825 3.325 143.100 3.555 ;
        RECT 141.105 1.260 141.335 2.390 ;
        RECT 141.825 1.490 142.055 3.325 ;
        RECT 143.345 2.920 143.575 4.350 ;
        RECT 142.310 2.690 143.575 2.920 ;
        RECT 143.345 1.260 143.575 2.390 ;
        RECT 144.065 2.300 144.295 4.080 ;
        RECT 144.525 3.250 145.040 4.230 ;
        RECT 145.405 4.015 145.635 4.580 ;
        RECT 146.150 3.280 146.775 4.305 ;
        RECT 147.425 3.785 147.655 4.580 ;
        RECT 144.525 2.690 145.410 3.250 ;
        RECT 145.790 2.300 146.075 3.050 ;
        RECT 144.065 2.065 146.075 2.300 ;
        RECT 144.065 1.490 144.450 2.065 ;
        RECT 145.350 1.260 145.690 1.750 ;
        RECT 146.305 1.500 146.775 3.280 ;
        RECT 147.425 3.325 148.700 3.555 ;
        RECT 147.425 1.490 147.655 3.325 ;
        RECT 148.945 2.920 149.175 4.350 ;
        RECT 149.665 3.785 149.895 4.580 ;
        RECT 147.910 2.690 149.175 2.920 ;
        RECT 149.665 3.325 150.940 3.555 ;
        RECT 148.945 1.260 149.175 2.390 ;
        RECT 149.665 1.490 149.895 3.325 ;
        RECT 151.185 2.920 151.415 4.350 ;
        RECT 151.905 3.785 152.135 4.580 ;
        RECT 150.150 2.690 151.415 2.920 ;
        RECT 151.905 3.325 153.180 3.555 ;
        RECT 151.185 1.260 151.415 2.390 ;
        RECT 151.905 1.490 152.135 3.325 ;
        RECT 153.425 2.920 153.655 4.350 ;
        RECT 154.290 3.695 154.630 4.580 ;
        RECT 155.265 3.785 155.495 4.580 ;
        RECT 155.265 3.325 156.540 3.555 ;
        RECT 152.390 2.690 153.655 2.920 ;
        RECT 153.425 1.260 153.655 2.390 ;
        RECT 154.290 1.260 154.630 2.950 ;
        RECT 155.265 1.490 155.495 3.325 ;
        RECT 156.785 2.920 157.015 4.350 ;
        RECT 157.505 3.785 157.735 4.580 ;
        RECT 155.750 2.690 157.015 2.920 ;
        RECT 157.505 3.325 158.780 3.555 ;
        RECT 156.785 1.260 157.015 2.390 ;
        RECT 157.505 1.490 157.735 3.325 ;
        RECT 159.025 2.920 159.255 4.350 ;
        RECT 159.745 3.785 159.975 4.580 ;
        RECT 157.990 2.690 159.255 2.920 ;
        RECT 159.745 3.325 161.020 3.555 ;
        RECT 159.025 1.260 159.255 2.390 ;
        RECT 159.745 1.490 159.975 3.325 ;
        RECT 161.265 2.920 161.495 4.350 ;
        RECT 161.985 3.785 162.215 4.580 ;
        RECT 160.230 2.690 161.495 2.920 ;
        RECT 161.985 3.325 163.260 3.555 ;
        RECT 161.265 1.260 161.495 2.390 ;
        RECT 161.985 1.490 162.215 3.325 ;
        RECT 163.505 2.920 163.735 4.350 ;
        RECT 164.225 3.785 164.455 4.580 ;
        RECT 162.470 2.690 163.735 2.920 ;
        RECT 164.225 3.325 165.500 3.555 ;
        RECT 163.505 1.260 163.735 2.390 ;
        RECT 164.225 1.490 164.455 3.325 ;
        RECT 165.745 2.920 165.975 4.350 ;
        RECT 164.710 2.690 165.975 2.920 ;
        RECT 165.745 1.260 165.975 2.390 ;
        RECT 166.465 2.300 166.695 4.080 ;
        RECT 166.925 3.250 167.440 4.230 ;
        RECT 167.805 4.015 168.035 4.580 ;
        RECT 168.550 3.280 169.175 4.305 ;
        RECT 169.825 3.785 170.055 4.580 ;
        RECT 166.925 2.690 167.810 3.250 ;
        RECT 168.190 2.300 168.475 3.050 ;
        RECT 166.465 2.065 168.475 2.300 ;
        RECT 166.465 1.490 166.850 2.065 ;
        RECT 167.750 1.260 168.090 1.750 ;
        RECT 168.705 1.500 169.175 3.280 ;
        RECT 169.825 3.325 171.100 3.555 ;
        RECT 169.825 1.490 170.055 3.325 ;
        RECT 171.345 2.920 171.575 4.350 ;
        RECT 172.065 3.785 172.295 4.580 ;
        RECT 170.310 2.690 171.575 2.920 ;
        RECT 172.065 3.325 173.340 3.555 ;
        RECT 171.345 1.260 171.575 2.390 ;
        RECT 172.065 1.490 172.295 3.325 ;
        RECT 173.585 2.920 173.815 4.350 ;
        RECT 174.430 3.690 174.770 4.580 ;
        RECT 172.550 2.690 173.815 2.920 ;
        RECT 173.585 1.260 173.815 2.390 ;
        RECT 174.430 1.260 174.770 2.960 ;
        RECT 57.170 0.660 175.180 1.260 ;
        RECT 57.170 0.610 57.550 0.660 ;
        RECT 57.900 0.620 58.340 0.660 ;
      LAYER Via1 ;
        RECT 2.190 59.990 2.450 60.250 ;
        RECT 20.035 59.990 20.295 60.250 ;
        RECT 0.825 58.805 1.085 59.065 ;
        RECT 0.825 58.145 1.085 58.405 ;
        RECT 0.825 57.485 1.085 57.745 ;
        RECT 0.825 56.825 1.085 57.085 ;
        RECT 0.825 56.165 1.085 56.425 ;
        RECT 0.825 55.505 1.085 55.765 ;
        RECT 0.825 54.845 1.085 55.105 ;
        RECT 0.825 54.185 1.085 54.445 ;
        RECT 0.825 53.525 1.085 53.785 ;
        RECT 0.825 52.865 1.085 53.125 ;
        RECT 0.825 52.205 1.085 52.465 ;
        RECT 0.825 51.545 1.085 51.805 ;
        RECT 0.825 50.885 1.085 51.145 ;
        RECT 0.825 50.225 1.085 50.485 ;
        RECT 5.310 47.865 5.570 48.125 ;
        RECT 5.970 47.865 6.230 48.125 ;
        RECT 6.630 47.865 6.890 48.125 ;
        RECT 5.310 47.205 5.570 47.465 ;
        RECT 5.970 47.205 6.230 47.465 ;
        RECT 6.630 47.205 6.890 47.465 ;
        RECT 5.310 46.545 5.570 46.805 ;
        RECT 5.970 46.545 6.230 46.805 ;
        RECT 6.630 46.545 6.890 46.805 ;
        RECT 5.310 22.265 5.570 22.525 ;
        RECT 5.970 22.265 6.230 22.525 ;
        RECT 6.630 22.265 6.890 22.525 ;
        RECT 5.310 21.605 5.570 21.865 ;
        RECT 5.970 21.605 6.230 21.865 ;
        RECT 6.630 21.605 6.890 21.865 ;
        RECT 5.310 20.945 5.570 21.205 ;
        RECT 5.970 20.945 6.230 21.205 ;
        RECT 6.630 20.945 6.890 21.205 ;
        RECT 11.115 58.805 11.375 59.065 ;
        RECT 11.115 58.145 11.375 58.405 ;
        RECT 11.115 57.485 11.375 57.745 ;
        RECT 11.115 56.825 11.375 57.085 ;
        RECT 11.115 56.165 11.375 56.425 ;
        RECT 11.115 55.505 11.375 55.765 ;
        RECT 11.115 54.845 11.375 55.105 ;
        RECT 11.115 54.185 11.375 54.445 ;
        RECT 11.115 53.525 11.375 53.785 ;
        RECT 11.115 52.865 11.375 53.125 ;
        RECT 11.115 52.205 11.375 52.465 ;
        RECT 11.115 51.545 11.375 51.805 ;
        RECT 11.115 50.885 11.375 51.145 ;
        RECT 11.115 50.225 11.375 50.485 ;
        RECT 24.185 59.990 24.445 60.250 ;
        RECT 42.030 59.990 42.290 60.250 ;
        RECT 15.610 45.165 15.870 45.425 ;
        RECT 16.270 45.165 16.530 45.425 ;
        RECT 16.930 45.165 17.190 45.425 ;
        RECT 15.610 44.505 15.870 44.765 ;
        RECT 16.270 44.505 16.530 44.765 ;
        RECT 16.930 44.505 17.190 44.765 ;
        RECT 15.610 43.845 15.870 44.105 ;
        RECT 16.270 43.845 16.530 44.105 ;
        RECT 16.930 43.845 17.190 44.105 ;
        RECT 15.610 24.965 15.870 25.225 ;
        RECT 16.270 24.965 16.530 25.225 ;
        RECT 16.930 24.965 17.190 25.225 ;
        RECT 15.610 24.305 15.870 24.565 ;
        RECT 16.270 24.305 16.530 24.565 ;
        RECT 16.930 24.305 17.190 24.565 ;
        RECT 15.610 23.645 15.870 23.905 ;
        RECT 16.270 23.645 16.530 23.905 ;
        RECT 16.930 23.645 17.190 23.905 ;
        RECT 9.750 8.805 10.010 9.065 ;
        RECT 21.400 58.805 21.660 59.065 ;
        RECT 21.400 58.145 21.660 58.405 ;
        RECT 21.400 57.485 21.660 57.745 ;
        RECT 21.400 56.825 21.660 57.085 ;
        RECT 21.400 56.165 21.660 56.425 ;
        RECT 21.400 55.505 21.660 55.765 ;
        RECT 21.400 54.845 21.660 55.105 ;
        RECT 21.400 54.185 21.660 54.445 ;
        RECT 21.400 53.525 21.660 53.785 ;
        RECT 21.400 52.865 21.660 53.125 ;
        RECT 21.400 52.205 21.660 52.465 ;
        RECT 21.400 51.545 21.660 51.805 ;
        RECT 21.400 50.885 21.660 51.145 ;
        RECT 21.400 50.225 21.660 50.485 ;
        RECT 22.820 58.805 23.080 59.065 ;
        RECT 22.820 58.145 23.080 58.405 ;
        RECT 22.820 57.485 23.080 57.745 ;
        RECT 22.820 56.825 23.080 57.085 ;
        RECT 22.820 56.165 23.080 56.425 ;
        RECT 22.820 55.505 23.080 55.765 ;
        RECT 22.820 54.845 23.080 55.105 ;
        RECT 22.820 54.185 23.080 54.445 ;
        RECT 22.820 53.525 23.080 53.785 ;
        RECT 22.820 52.865 23.080 53.125 ;
        RECT 22.820 52.205 23.080 52.465 ;
        RECT 22.820 51.545 23.080 51.805 ;
        RECT 22.820 50.885 23.080 51.145 ;
        RECT 22.820 50.225 23.080 50.485 ;
        RECT 27.305 47.865 27.565 48.125 ;
        RECT 27.965 47.865 28.225 48.125 ;
        RECT 28.625 47.865 28.885 48.125 ;
        RECT 27.305 47.205 27.565 47.465 ;
        RECT 27.965 47.205 28.225 47.465 ;
        RECT 28.625 47.205 28.885 47.465 ;
        RECT 27.305 46.545 27.565 46.805 ;
        RECT 27.965 46.545 28.225 46.805 ;
        RECT 28.625 46.545 28.885 46.805 ;
        RECT 27.305 22.265 27.565 22.525 ;
        RECT 27.965 22.265 28.225 22.525 ;
        RECT 28.625 22.265 28.885 22.525 ;
        RECT 27.305 21.605 27.565 21.865 ;
        RECT 27.965 21.605 28.225 21.865 ;
        RECT 28.625 21.605 28.885 21.865 ;
        RECT 27.305 20.945 27.565 21.205 ;
        RECT 27.965 20.945 28.225 21.205 ;
        RECT 28.625 20.945 28.885 21.205 ;
        RECT 33.110 58.805 33.370 59.065 ;
        RECT 33.110 58.145 33.370 58.405 ;
        RECT 33.110 57.485 33.370 57.745 ;
        RECT 33.110 56.825 33.370 57.085 ;
        RECT 33.110 56.165 33.370 56.425 ;
        RECT 33.110 55.505 33.370 55.765 ;
        RECT 33.110 54.845 33.370 55.105 ;
        RECT 33.110 54.185 33.370 54.445 ;
        RECT 33.110 53.525 33.370 53.785 ;
        RECT 33.110 52.865 33.370 53.125 ;
        RECT 33.110 52.205 33.370 52.465 ;
        RECT 33.110 51.545 33.370 51.805 ;
        RECT 33.110 50.885 33.370 51.145 ;
        RECT 33.110 50.225 33.370 50.485 ;
        RECT 46.180 59.990 46.440 60.250 ;
        RECT 64.025 59.990 64.285 60.250 ;
        RECT 37.605 45.165 37.865 45.425 ;
        RECT 38.265 45.165 38.525 45.425 ;
        RECT 38.925 45.165 39.185 45.425 ;
        RECT 37.605 44.505 37.865 44.765 ;
        RECT 38.265 44.505 38.525 44.765 ;
        RECT 38.925 44.505 39.185 44.765 ;
        RECT 37.605 43.845 37.865 44.105 ;
        RECT 38.265 43.845 38.525 44.105 ;
        RECT 38.925 43.845 39.185 44.105 ;
        RECT 37.605 24.965 37.865 25.225 ;
        RECT 38.265 24.965 38.525 25.225 ;
        RECT 38.925 24.965 39.185 25.225 ;
        RECT 37.605 24.305 37.865 24.565 ;
        RECT 38.265 24.305 38.525 24.565 ;
        RECT 38.925 24.305 39.185 24.565 ;
        RECT 37.605 23.645 37.865 23.905 ;
        RECT 38.265 23.645 38.525 23.905 ;
        RECT 38.925 23.645 39.185 23.905 ;
        RECT 12.480 8.805 12.740 9.065 ;
        RECT 31.745 8.805 32.005 9.065 ;
        RECT 43.395 58.805 43.655 59.065 ;
        RECT 43.395 58.145 43.655 58.405 ;
        RECT 43.395 57.485 43.655 57.745 ;
        RECT 43.395 56.825 43.655 57.085 ;
        RECT 43.395 56.165 43.655 56.425 ;
        RECT 43.395 55.505 43.655 55.765 ;
        RECT 43.395 54.845 43.655 55.105 ;
        RECT 43.395 54.185 43.655 54.445 ;
        RECT 43.395 53.525 43.655 53.785 ;
        RECT 43.395 52.865 43.655 53.125 ;
        RECT 43.395 52.205 43.655 52.465 ;
        RECT 43.395 51.545 43.655 51.805 ;
        RECT 43.395 50.885 43.655 51.145 ;
        RECT 43.395 50.225 43.655 50.485 ;
        RECT 44.815 58.805 45.075 59.065 ;
        RECT 44.815 58.145 45.075 58.405 ;
        RECT 44.815 57.485 45.075 57.745 ;
        RECT 44.815 56.825 45.075 57.085 ;
        RECT 44.815 56.165 45.075 56.425 ;
        RECT 44.815 55.505 45.075 55.765 ;
        RECT 44.815 54.845 45.075 55.105 ;
        RECT 44.815 54.185 45.075 54.445 ;
        RECT 44.815 53.525 45.075 53.785 ;
        RECT 44.815 52.865 45.075 53.125 ;
        RECT 44.815 52.205 45.075 52.465 ;
        RECT 44.815 51.545 45.075 51.805 ;
        RECT 44.815 50.885 45.075 51.145 ;
        RECT 44.815 50.225 45.075 50.485 ;
        RECT 49.300 47.865 49.560 48.125 ;
        RECT 49.960 47.865 50.220 48.125 ;
        RECT 50.620 47.865 50.880 48.125 ;
        RECT 49.300 47.205 49.560 47.465 ;
        RECT 49.960 47.205 50.220 47.465 ;
        RECT 50.620 47.205 50.880 47.465 ;
        RECT 49.300 46.545 49.560 46.805 ;
        RECT 49.960 46.545 50.220 46.805 ;
        RECT 50.620 46.545 50.880 46.805 ;
        RECT 49.300 22.265 49.560 22.525 ;
        RECT 49.960 22.265 50.220 22.525 ;
        RECT 50.620 22.265 50.880 22.525 ;
        RECT 49.300 21.605 49.560 21.865 ;
        RECT 49.960 21.605 50.220 21.865 ;
        RECT 50.620 21.605 50.880 21.865 ;
        RECT 49.300 20.945 49.560 21.205 ;
        RECT 49.960 20.945 50.220 21.205 ;
        RECT 50.620 20.945 50.880 21.205 ;
        RECT 55.105 58.805 55.365 59.065 ;
        RECT 55.105 58.145 55.365 58.405 ;
        RECT 55.105 57.485 55.365 57.745 ;
        RECT 55.105 56.825 55.365 57.085 ;
        RECT 55.105 56.165 55.365 56.425 ;
        RECT 55.105 55.505 55.365 55.765 ;
        RECT 55.105 54.845 55.365 55.105 ;
        RECT 55.105 54.185 55.365 54.445 ;
        RECT 55.105 53.525 55.365 53.785 ;
        RECT 55.105 52.865 55.365 53.125 ;
        RECT 55.105 52.205 55.365 52.465 ;
        RECT 55.105 51.545 55.365 51.805 ;
        RECT 55.105 50.885 55.365 51.145 ;
        RECT 55.105 50.225 55.365 50.485 ;
        RECT 68.175 59.990 68.435 60.250 ;
        RECT 86.020 59.990 86.280 60.250 ;
        RECT 59.600 45.165 59.860 45.425 ;
        RECT 60.260 45.165 60.520 45.425 ;
        RECT 60.920 45.165 61.180 45.425 ;
        RECT 59.600 44.505 59.860 44.765 ;
        RECT 60.260 44.505 60.520 44.765 ;
        RECT 60.920 44.505 61.180 44.765 ;
        RECT 59.600 43.845 59.860 44.105 ;
        RECT 60.260 43.845 60.520 44.105 ;
        RECT 60.920 43.845 61.180 44.105 ;
        RECT 59.600 24.965 59.860 25.225 ;
        RECT 60.260 24.965 60.520 25.225 ;
        RECT 60.920 24.965 61.180 25.225 ;
        RECT 59.600 24.305 59.860 24.565 ;
        RECT 60.260 24.305 60.520 24.565 ;
        RECT 60.920 24.305 61.180 24.565 ;
        RECT 59.600 23.645 59.860 23.905 ;
        RECT 60.260 23.645 60.520 23.905 ;
        RECT 60.920 23.645 61.180 23.905 ;
        RECT 34.475 8.805 34.735 9.065 ;
        RECT 53.740 8.805 54.000 9.065 ;
        RECT 65.390 58.805 65.650 59.065 ;
        RECT 65.390 58.145 65.650 58.405 ;
        RECT 65.390 57.485 65.650 57.745 ;
        RECT 65.390 56.825 65.650 57.085 ;
        RECT 65.390 56.165 65.650 56.425 ;
        RECT 65.390 55.505 65.650 55.765 ;
        RECT 65.390 54.845 65.650 55.105 ;
        RECT 65.390 54.185 65.650 54.445 ;
        RECT 65.390 53.525 65.650 53.785 ;
        RECT 65.390 52.865 65.650 53.125 ;
        RECT 65.390 52.205 65.650 52.465 ;
        RECT 65.390 51.545 65.650 51.805 ;
        RECT 65.390 50.885 65.650 51.145 ;
        RECT 65.390 50.225 65.650 50.485 ;
        RECT 66.810 58.805 67.070 59.065 ;
        RECT 66.810 58.145 67.070 58.405 ;
        RECT 66.810 57.485 67.070 57.745 ;
        RECT 66.810 56.825 67.070 57.085 ;
        RECT 66.810 56.165 67.070 56.425 ;
        RECT 66.810 55.505 67.070 55.765 ;
        RECT 66.810 54.845 67.070 55.105 ;
        RECT 66.810 54.185 67.070 54.445 ;
        RECT 66.810 53.525 67.070 53.785 ;
        RECT 66.810 52.865 67.070 53.125 ;
        RECT 66.810 52.205 67.070 52.465 ;
        RECT 66.810 51.545 67.070 51.805 ;
        RECT 66.810 50.885 67.070 51.145 ;
        RECT 66.810 50.225 67.070 50.485 ;
        RECT 71.295 47.865 71.555 48.125 ;
        RECT 71.955 47.865 72.215 48.125 ;
        RECT 72.615 47.865 72.875 48.125 ;
        RECT 71.295 47.205 71.555 47.465 ;
        RECT 71.955 47.205 72.215 47.465 ;
        RECT 72.615 47.205 72.875 47.465 ;
        RECT 71.295 46.545 71.555 46.805 ;
        RECT 71.955 46.545 72.215 46.805 ;
        RECT 72.615 46.545 72.875 46.805 ;
        RECT 71.295 22.265 71.555 22.525 ;
        RECT 71.955 22.265 72.215 22.525 ;
        RECT 72.615 22.265 72.875 22.525 ;
        RECT 71.295 21.605 71.555 21.865 ;
        RECT 71.955 21.605 72.215 21.865 ;
        RECT 72.615 21.605 72.875 21.865 ;
        RECT 71.295 20.945 71.555 21.205 ;
        RECT 71.955 20.945 72.215 21.205 ;
        RECT 72.615 20.945 72.875 21.205 ;
        RECT 77.100 58.805 77.360 59.065 ;
        RECT 77.100 58.145 77.360 58.405 ;
        RECT 77.100 57.485 77.360 57.745 ;
        RECT 77.100 56.825 77.360 57.085 ;
        RECT 77.100 56.165 77.360 56.425 ;
        RECT 77.100 55.505 77.360 55.765 ;
        RECT 77.100 54.845 77.360 55.105 ;
        RECT 77.100 54.185 77.360 54.445 ;
        RECT 77.100 53.525 77.360 53.785 ;
        RECT 77.100 52.865 77.360 53.125 ;
        RECT 77.100 52.205 77.360 52.465 ;
        RECT 77.100 51.545 77.360 51.805 ;
        RECT 77.100 50.885 77.360 51.145 ;
        RECT 77.100 50.225 77.360 50.485 ;
        RECT 90.170 59.990 90.430 60.250 ;
        RECT 108.015 59.990 108.275 60.250 ;
        RECT 81.595 45.165 81.855 45.425 ;
        RECT 82.255 45.165 82.515 45.425 ;
        RECT 82.915 45.165 83.175 45.425 ;
        RECT 81.595 44.505 81.855 44.765 ;
        RECT 82.255 44.505 82.515 44.765 ;
        RECT 82.915 44.505 83.175 44.765 ;
        RECT 81.595 43.845 81.855 44.105 ;
        RECT 82.255 43.845 82.515 44.105 ;
        RECT 82.915 43.845 83.175 44.105 ;
        RECT 81.595 24.965 81.855 25.225 ;
        RECT 82.255 24.965 82.515 25.225 ;
        RECT 82.915 24.965 83.175 25.225 ;
        RECT 81.595 24.305 81.855 24.565 ;
        RECT 82.255 24.305 82.515 24.565 ;
        RECT 82.915 24.305 83.175 24.565 ;
        RECT 81.595 23.645 81.855 23.905 ;
        RECT 82.255 23.645 82.515 23.905 ;
        RECT 82.915 23.645 83.175 23.905 ;
        RECT 56.470 8.805 56.730 9.065 ;
        RECT 75.735 8.805 75.995 9.065 ;
        RECT 87.385 58.805 87.645 59.065 ;
        RECT 87.385 58.145 87.645 58.405 ;
        RECT 87.385 57.485 87.645 57.745 ;
        RECT 87.385 56.825 87.645 57.085 ;
        RECT 87.385 56.165 87.645 56.425 ;
        RECT 87.385 55.505 87.645 55.765 ;
        RECT 87.385 54.845 87.645 55.105 ;
        RECT 87.385 54.185 87.645 54.445 ;
        RECT 87.385 53.525 87.645 53.785 ;
        RECT 87.385 52.865 87.645 53.125 ;
        RECT 87.385 52.205 87.645 52.465 ;
        RECT 87.385 51.545 87.645 51.805 ;
        RECT 87.385 50.885 87.645 51.145 ;
        RECT 87.385 50.225 87.645 50.485 ;
        RECT 88.805 58.805 89.065 59.065 ;
        RECT 88.805 58.145 89.065 58.405 ;
        RECT 88.805 57.485 89.065 57.745 ;
        RECT 88.805 56.825 89.065 57.085 ;
        RECT 88.805 56.165 89.065 56.425 ;
        RECT 88.805 55.505 89.065 55.765 ;
        RECT 88.805 54.845 89.065 55.105 ;
        RECT 88.805 54.185 89.065 54.445 ;
        RECT 88.805 53.525 89.065 53.785 ;
        RECT 88.805 52.865 89.065 53.125 ;
        RECT 88.805 52.205 89.065 52.465 ;
        RECT 88.805 51.545 89.065 51.805 ;
        RECT 88.805 50.885 89.065 51.145 ;
        RECT 88.805 50.225 89.065 50.485 ;
        RECT 93.290 47.865 93.550 48.125 ;
        RECT 93.950 47.865 94.210 48.125 ;
        RECT 94.610 47.865 94.870 48.125 ;
        RECT 93.290 47.205 93.550 47.465 ;
        RECT 93.950 47.205 94.210 47.465 ;
        RECT 94.610 47.205 94.870 47.465 ;
        RECT 93.290 46.545 93.550 46.805 ;
        RECT 93.950 46.545 94.210 46.805 ;
        RECT 94.610 46.545 94.870 46.805 ;
        RECT 93.290 22.265 93.550 22.525 ;
        RECT 93.950 22.265 94.210 22.525 ;
        RECT 94.610 22.265 94.870 22.525 ;
        RECT 93.290 21.605 93.550 21.865 ;
        RECT 93.950 21.605 94.210 21.865 ;
        RECT 94.610 21.605 94.870 21.865 ;
        RECT 93.290 20.945 93.550 21.205 ;
        RECT 93.950 20.945 94.210 21.205 ;
        RECT 94.610 20.945 94.870 21.205 ;
        RECT 99.095 58.805 99.355 59.065 ;
        RECT 99.095 58.145 99.355 58.405 ;
        RECT 99.095 57.485 99.355 57.745 ;
        RECT 99.095 56.825 99.355 57.085 ;
        RECT 99.095 56.165 99.355 56.425 ;
        RECT 99.095 55.505 99.355 55.765 ;
        RECT 99.095 54.845 99.355 55.105 ;
        RECT 99.095 54.185 99.355 54.445 ;
        RECT 99.095 53.525 99.355 53.785 ;
        RECT 99.095 52.865 99.355 53.125 ;
        RECT 99.095 52.205 99.355 52.465 ;
        RECT 99.095 51.545 99.355 51.805 ;
        RECT 99.095 50.885 99.355 51.145 ;
        RECT 99.095 50.225 99.355 50.485 ;
        RECT 112.165 59.990 112.425 60.250 ;
        RECT 130.010 59.990 130.270 60.250 ;
        RECT 103.590 45.165 103.850 45.425 ;
        RECT 104.250 45.165 104.510 45.425 ;
        RECT 104.910 45.165 105.170 45.425 ;
        RECT 103.590 44.505 103.850 44.765 ;
        RECT 104.250 44.505 104.510 44.765 ;
        RECT 104.910 44.505 105.170 44.765 ;
        RECT 103.590 43.845 103.850 44.105 ;
        RECT 104.250 43.845 104.510 44.105 ;
        RECT 104.910 43.845 105.170 44.105 ;
        RECT 103.590 24.965 103.850 25.225 ;
        RECT 104.250 24.965 104.510 25.225 ;
        RECT 104.910 24.965 105.170 25.225 ;
        RECT 103.590 24.305 103.850 24.565 ;
        RECT 104.250 24.305 104.510 24.565 ;
        RECT 104.910 24.305 105.170 24.565 ;
        RECT 103.590 23.645 103.850 23.905 ;
        RECT 104.250 23.645 104.510 23.905 ;
        RECT 104.910 23.645 105.170 23.905 ;
        RECT 78.465 8.805 78.725 9.065 ;
        RECT 97.730 8.805 97.990 9.065 ;
        RECT 109.380 58.805 109.640 59.065 ;
        RECT 109.380 58.145 109.640 58.405 ;
        RECT 109.380 57.485 109.640 57.745 ;
        RECT 109.380 56.825 109.640 57.085 ;
        RECT 109.380 56.165 109.640 56.425 ;
        RECT 109.380 55.505 109.640 55.765 ;
        RECT 109.380 54.845 109.640 55.105 ;
        RECT 109.380 54.185 109.640 54.445 ;
        RECT 109.380 53.525 109.640 53.785 ;
        RECT 109.380 52.865 109.640 53.125 ;
        RECT 109.380 52.205 109.640 52.465 ;
        RECT 109.380 51.545 109.640 51.805 ;
        RECT 109.380 50.885 109.640 51.145 ;
        RECT 109.380 50.225 109.640 50.485 ;
        RECT 110.800 58.805 111.060 59.065 ;
        RECT 110.800 58.145 111.060 58.405 ;
        RECT 110.800 57.485 111.060 57.745 ;
        RECT 110.800 56.825 111.060 57.085 ;
        RECT 110.800 56.165 111.060 56.425 ;
        RECT 110.800 55.505 111.060 55.765 ;
        RECT 110.800 54.845 111.060 55.105 ;
        RECT 110.800 54.185 111.060 54.445 ;
        RECT 110.800 53.525 111.060 53.785 ;
        RECT 110.800 52.865 111.060 53.125 ;
        RECT 110.800 52.205 111.060 52.465 ;
        RECT 110.800 51.545 111.060 51.805 ;
        RECT 110.800 50.885 111.060 51.145 ;
        RECT 110.800 50.225 111.060 50.485 ;
        RECT 115.285 47.865 115.545 48.125 ;
        RECT 115.945 47.865 116.205 48.125 ;
        RECT 116.605 47.865 116.865 48.125 ;
        RECT 115.285 47.205 115.545 47.465 ;
        RECT 115.945 47.205 116.205 47.465 ;
        RECT 116.605 47.205 116.865 47.465 ;
        RECT 115.285 46.545 115.545 46.805 ;
        RECT 115.945 46.545 116.205 46.805 ;
        RECT 116.605 46.545 116.865 46.805 ;
        RECT 115.285 22.265 115.545 22.525 ;
        RECT 115.945 22.265 116.205 22.525 ;
        RECT 116.605 22.265 116.865 22.525 ;
        RECT 115.285 21.605 115.545 21.865 ;
        RECT 115.945 21.605 116.205 21.865 ;
        RECT 116.605 21.605 116.865 21.865 ;
        RECT 115.285 20.945 115.545 21.205 ;
        RECT 115.945 20.945 116.205 21.205 ;
        RECT 116.605 20.945 116.865 21.205 ;
        RECT 121.090 58.805 121.350 59.065 ;
        RECT 121.090 58.145 121.350 58.405 ;
        RECT 121.090 57.485 121.350 57.745 ;
        RECT 121.090 56.825 121.350 57.085 ;
        RECT 121.090 56.165 121.350 56.425 ;
        RECT 121.090 55.505 121.350 55.765 ;
        RECT 121.090 54.845 121.350 55.105 ;
        RECT 121.090 54.185 121.350 54.445 ;
        RECT 121.090 53.525 121.350 53.785 ;
        RECT 121.090 52.865 121.350 53.125 ;
        RECT 121.090 52.205 121.350 52.465 ;
        RECT 121.090 51.545 121.350 51.805 ;
        RECT 121.090 50.885 121.350 51.145 ;
        RECT 121.090 50.225 121.350 50.485 ;
        RECT 134.160 59.990 134.420 60.250 ;
        RECT 152.005 59.990 152.265 60.250 ;
        RECT 125.585 45.165 125.845 45.425 ;
        RECT 126.245 45.165 126.505 45.425 ;
        RECT 126.905 45.165 127.165 45.425 ;
        RECT 125.585 44.505 125.845 44.765 ;
        RECT 126.245 44.505 126.505 44.765 ;
        RECT 126.905 44.505 127.165 44.765 ;
        RECT 125.585 43.845 125.845 44.105 ;
        RECT 126.245 43.845 126.505 44.105 ;
        RECT 126.905 43.845 127.165 44.105 ;
        RECT 125.585 24.965 125.845 25.225 ;
        RECT 126.245 24.965 126.505 25.225 ;
        RECT 126.905 24.965 127.165 25.225 ;
        RECT 125.585 24.305 125.845 24.565 ;
        RECT 126.245 24.305 126.505 24.565 ;
        RECT 126.905 24.305 127.165 24.565 ;
        RECT 125.585 23.645 125.845 23.905 ;
        RECT 126.245 23.645 126.505 23.905 ;
        RECT 126.905 23.645 127.165 23.905 ;
        RECT 100.460 8.805 100.720 9.065 ;
        RECT 119.725 8.805 119.985 9.065 ;
        RECT 131.375 58.805 131.635 59.065 ;
        RECT 131.375 58.145 131.635 58.405 ;
        RECT 131.375 57.485 131.635 57.745 ;
        RECT 131.375 56.825 131.635 57.085 ;
        RECT 131.375 56.165 131.635 56.425 ;
        RECT 131.375 55.505 131.635 55.765 ;
        RECT 131.375 54.845 131.635 55.105 ;
        RECT 131.375 54.185 131.635 54.445 ;
        RECT 131.375 53.525 131.635 53.785 ;
        RECT 131.375 52.865 131.635 53.125 ;
        RECT 131.375 52.205 131.635 52.465 ;
        RECT 131.375 51.545 131.635 51.805 ;
        RECT 131.375 50.885 131.635 51.145 ;
        RECT 131.375 50.225 131.635 50.485 ;
        RECT 132.795 58.805 133.055 59.065 ;
        RECT 132.795 58.145 133.055 58.405 ;
        RECT 132.795 57.485 133.055 57.745 ;
        RECT 132.795 56.825 133.055 57.085 ;
        RECT 132.795 56.165 133.055 56.425 ;
        RECT 132.795 55.505 133.055 55.765 ;
        RECT 132.795 54.845 133.055 55.105 ;
        RECT 132.795 54.185 133.055 54.445 ;
        RECT 132.795 53.525 133.055 53.785 ;
        RECT 132.795 52.865 133.055 53.125 ;
        RECT 132.795 52.205 133.055 52.465 ;
        RECT 132.795 51.545 133.055 51.805 ;
        RECT 132.795 50.885 133.055 51.145 ;
        RECT 132.795 50.225 133.055 50.485 ;
        RECT 137.280 47.865 137.540 48.125 ;
        RECT 137.940 47.865 138.200 48.125 ;
        RECT 138.600 47.865 138.860 48.125 ;
        RECT 137.280 47.205 137.540 47.465 ;
        RECT 137.940 47.205 138.200 47.465 ;
        RECT 138.600 47.205 138.860 47.465 ;
        RECT 137.280 46.545 137.540 46.805 ;
        RECT 137.940 46.545 138.200 46.805 ;
        RECT 138.600 46.545 138.860 46.805 ;
        RECT 137.280 22.265 137.540 22.525 ;
        RECT 137.940 22.265 138.200 22.525 ;
        RECT 138.600 22.265 138.860 22.525 ;
        RECT 137.280 21.605 137.540 21.865 ;
        RECT 137.940 21.605 138.200 21.865 ;
        RECT 138.600 21.605 138.860 21.865 ;
        RECT 137.280 20.945 137.540 21.205 ;
        RECT 137.940 20.945 138.200 21.205 ;
        RECT 138.600 20.945 138.860 21.205 ;
        RECT 143.085 58.805 143.345 59.065 ;
        RECT 143.085 58.145 143.345 58.405 ;
        RECT 143.085 57.485 143.345 57.745 ;
        RECT 143.085 56.825 143.345 57.085 ;
        RECT 143.085 56.165 143.345 56.425 ;
        RECT 143.085 55.505 143.345 55.765 ;
        RECT 143.085 54.845 143.345 55.105 ;
        RECT 143.085 54.185 143.345 54.445 ;
        RECT 143.085 53.525 143.345 53.785 ;
        RECT 143.085 52.865 143.345 53.125 ;
        RECT 143.085 52.205 143.345 52.465 ;
        RECT 143.085 51.545 143.345 51.805 ;
        RECT 143.085 50.885 143.345 51.145 ;
        RECT 143.085 50.225 143.345 50.485 ;
        RECT 156.155 59.990 156.415 60.250 ;
        RECT 174.000 59.990 174.260 60.250 ;
        RECT 147.580 45.165 147.840 45.425 ;
        RECT 148.240 45.165 148.500 45.425 ;
        RECT 148.900 45.165 149.160 45.425 ;
        RECT 147.580 44.505 147.840 44.765 ;
        RECT 148.240 44.505 148.500 44.765 ;
        RECT 148.900 44.505 149.160 44.765 ;
        RECT 147.580 43.845 147.840 44.105 ;
        RECT 148.240 43.845 148.500 44.105 ;
        RECT 148.900 43.845 149.160 44.105 ;
        RECT 147.580 24.965 147.840 25.225 ;
        RECT 148.240 24.965 148.500 25.225 ;
        RECT 148.900 24.965 149.160 25.225 ;
        RECT 147.580 24.305 147.840 24.565 ;
        RECT 148.240 24.305 148.500 24.565 ;
        RECT 148.900 24.305 149.160 24.565 ;
        RECT 147.580 23.645 147.840 23.905 ;
        RECT 148.240 23.645 148.500 23.905 ;
        RECT 148.900 23.645 149.160 23.905 ;
        RECT 122.455 8.805 122.715 9.065 ;
        RECT 141.720 8.805 141.980 9.065 ;
        RECT 153.370 58.805 153.630 59.065 ;
        RECT 153.370 58.145 153.630 58.405 ;
        RECT 153.370 57.485 153.630 57.745 ;
        RECT 153.370 56.825 153.630 57.085 ;
        RECT 153.370 56.165 153.630 56.425 ;
        RECT 153.370 55.505 153.630 55.765 ;
        RECT 153.370 54.845 153.630 55.105 ;
        RECT 153.370 54.185 153.630 54.445 ;
        RECT 153.370 53.525 153.630 53.785 ;
        RECT 153.370 52.865 153.630 53.125 ;
        RECT 153.370 52.205 153.630 52.465 ;
        RECT 153.370 51.545 153.630 51.805 ;
        RECT 153.370 50.885 153.630 51.145 ;
        RECT 153.370 50.225 153.630 50.485 ;
        RECT 154.790 58.805 155.050 59.065 ;
        RECT 154.790 58.145 155.050 58.405 ;
        RECT 154.790 57.485 155.050 57.745 ;
        RECT 154.790 56.825 155.050 57.085 ;
        RECT 154.790 56.165 155.050 56.425 ;
        RECT 154.790 55.505 155.050 55.765 ;
        RECT 154.790 54.845 155.050 55.105 ;
        RECT 154.790 54.185 155.050 54.445 ;
        RECT 154.790 53.525 155.050 53.785 ;
        RECT 154.790 52.865 155.050 53.125 ;
        RECT 154.790 52.205 155.050 52.465 ;
        RECT 154.790 51.545 155.050 51.805 ;
        RECT 154.790 50.885 155.050 51.145 ;
        RECT 154.790 50.225 155.050 50.485 ;
        RECT 159.275 47.865 159.535 48.125 ;
        RECT 159.935 47.865 160.195 48.125 ;
        RECT 160.595 47.865 160.855 48.125 ;
        RECT 159.275 47.205 159.535 47.465 ;
        RECT 159.935 47.205 160.195 47.465 ;
        RECT 160.595 47.205 160.855 47.465 ;
        RECT 159.275 46.545 159.535 46.805 ;
        RECT 159.935 46.545 160.195 46.805 ;
        RECT 160.595 46.545 160.855 46.805 ;
        RECT 159.275 22.265 159.535 22.525 ;
        RECT 159.935 22.265 160.195 22.525 ;
        RECT 160.595 22.265 160.855 22.525 ;
        RECT 159.275 21.605 159.535 21.865 ;
        RECT 159.935 21.605 160.195 21.865 ;
        RECT 160.595 21.605 160.855 21.865 ;
        RECT 159.275 20.945 159.535 21.205 ;
        RECT 159.935 20.945 160.195 21.205 ;
        RECT 160.595 20.945 160.855 21.205 ;
        RECT 165.080 58.805 165.340 59.065 ;
        RECT 165.080 58.145 165.340 58.405 ;
        RECT 165.080 57.485 165.340 57.745 ;
        RECT 165.080 56.825 165.340 57.085 ;
        RECT 165.080 56.165 165.340 56.425 ;
        RECT 165.080 55.505 165.340 55.765 ;
        RECT 165.080 54.845 165.340 55.105 ;
        RECT 165.080 54.185 165.340 54.445 ;
        RECT 165.080 53.525 165.340 53.785 ;
        RECT 165.080 52.865 165.340 53.125 ;
        RECT 165.080 52.205 165.340 52.465 ;
        RECT 165.080 51.545 165.340 51.805 ;
        RECT 165.080 50.885 165.340 51.145 ;
        RECT 165.080 50.225 165.340 50.485 ;
        RECT 169.575 45.165 169.835 45.425 ;
        RECT 170.235 45.165 170.495 45.425 ;
        RECT 170.895 45.165 171.155 45.425 ;
        RECT 169.575 44.505 169.835 44.765 ;
        RECT 170.235 44.505 170.495 44.765 ;
        RECT 170.895 44.505 171.155 44.765 ;
        RECT 169.575 43.845 169.835 44.105 ;
        RECT 170.235 43.845 170.495 44.105 ;
        RECT 170.895 43.845 171.155 44.105 ;
        RECT 169.575 24.965 169.835 25.225 ;
        RECT 170.235 24.965 170.495 25.225 ;
        RECT 170.895 24.965 171.155 25.225 ;
        RECT 169.575 24.305 169.835 24.565 ;
        RECT 170.235 24.305 170.495 24.565 ;
        RECT 170.895 24.305 171.155 24.565 ;
        RECT 169.575 23.645 169.835 23.905 ;
        RECT 170.235 23.645 170.495 23.905 ;
        RECT 170.895 23.645 171.155 23.905 ;
        RECT 144.450 8.805 144.710 9.065 ;
        RECT 163.715 8.805 163.975 9.065 ;
        RECT 175.365 58.805 175.625 59.065 ;
        RECT 175.365 58.145 175.625 58.405 ;
        RECT 175.365 57.485 175.625 57.745 ;
        RECT 175.365 56.825 175.625 57.085 ;
        RECT 175.365 56.165 175.625 56.425 ;
        RECT 175.365 55.505 175.625 55.765 ;
        RECT 175.365 54.845 175.625 55.105 ;
        RECT 175.365 54.185 175.625 54.445 ;
        RECT 175.365 53.525 175.625 53.785 ;
        RECT 175.365 52.865 175.625 53.125 ;
        RECT 175.365 52.205 175.625 52.465 ;
        RECT 175.365 51.545 175.625 51.805 ;
        RECT 175.365 50.885 175.625 51.145 ;
        RECT 175.365 50.225 175.625 50.485 ;
        RECT 177.210 55.175 177.470 55.435 ;
        RECT 177.210 54.515 177.470 54.775 ;
        RECT 177.210 53.855 177.470 54.115 ;
        RECT 177.210 53.195 177.470 53.455 ;
        RECT 177.210 52.535 177.470 52.795 ;
        RECT 177.210 51.875 177.470 52.135 ;
        RECT 177.210 51.215 177.470 51.475 ;
        RECT 177.210 50.555 177.470 50.815 ;
        RECT 177.210 18.175 177.470 18.435 ;
        RECT 177.210 17.515 177.470 17.775 ;
        RECT 177.210 16.855 177.470 17.115 ;
        RECT 177.210 16.195 177.470 16.455 ;
        RECT 177.210 15.535 177.470 15.795 ;
        RECT 177.210 14.875 177.470 15.135 ;
        RECT 177.210 14.215 177.470 14.475 ;
        RECT 177.210 13.555 177.470 13.815 ;
        RECT 177.210 12.895 177.470 13.155 ;
        RECT 177.210 12.235 177.470 12.495 ;
        RECT 177.210 11.575 177.470 11.835 ;
        RECT 177.210 10.915 177.470 11.175 ;
        RECT 177.210 10.255 177.470 10.515 ;
        RECT 177.210 9.595 177.470 9.855 ;
        RECT 166.445 8.805 166.705 9.065 ;
        RECT 177.210 8.935 177.470 9.195 ;
        RECT 178.995 55.175 179.255 55.435 ;
        RECT 181.850 55.175 182.110 55.435 ;
        RECT 178.995 54.515 179.255 54.775 ;
        RECT 181.850 54.515 182.110 54.775 ;
        RECT 178.995 53.855 179.255 54.115 ;
        RECT 181.850 53.855 182.110 54.115 ;
        RECT 178.995 53.195 179.255 53.455 ;
        RECT 181.850 53.195 182.110 53.455 ;
        RECT 178.995 52.535 179.255 52.795 ;
        RECT 181.850 52.535 182.110 52.795 ;
        RECT 178.995 51.875 179.255 52.135 ;
        RECT 181.850 51.875 182.110 52.135 ;
        RECT 178.995 51.215 179.255 51.475 ;
        RECT 181.850 51.215 182.110 51.475 ;
        RECT 178.995 50.555 179.255 50.815 ;
        RECT 181.850 50.555 182.110 50.815 ;
        RECT 177.970 47.865 178.230 48.125 ;
        RECT 177.970 47.205 178.230 47.465 ;
        RECT 177.970 46.545 178.230 46.805 ;
        RECT 178.995 18.175 179.255 18.435 ;
        RECT 181.850 18.175 182.110 18.435 ;
        RECT 178.995 17.515 179.255 17.775 ;
        RECT 181.850 17.515 182.110 17.775 ;
        RECT 178.995 16.855 179.255 17.115 ;
        RECT 181.850 16.855 182.110 17.115 ;
        RECT 178.995 16.195 179.255 16.455 ;
        RECT 181.850 16.195 182.110 16.455 ;
        RECT 178.995 15.535 179.255 15.795 ;
        RECT 181.850 15.535 182.110 15.795 ;
        RECT 178.995 14.875 179.255 15.135 ;
        RECT 181.850 14.875 182.110 15.135 ;
        RECT 178.995 14.215 179.255 14.475 ;
        RECT 181.850 14.215 182.110 14.475 ;
        RECT 178.995 13.555 179.255 13.815 ;
        RECT 181.850 13.555 182.110 13.815 ;
        RECT 178.995 12.895 179.255 13.155 ;
        RECT 181.850 12.895 182.110 13.155 ;
        RECT 178.995 12.235 179.255 12.495 ;
        RECT 181.850 12.235 182.110 12.495 ;
        RECT 178.995 11.575 179.255 11.835 ;
        RECT 181.850 11.575 182.110 11.835 ;
        RECT 178.995 10.915 179.255 11.175 ;
        RECT 181.850 10.915 182.110 11.175 ;
        RECT 178.995 10.255 179.255 10.515 ;
        RECT 181.850 10.255 182.110 10.515 ;
        RECT 178.995 9.595 179.255 9.855 ;
        RECT 181.850 9.595 182.110 9.855 ;
        RECT 178.995 8.935 179.255 9.195 ;
        RECT 181.850 8.935 182.110 9.195 ;
        RECT 183.635 55.175 183.895 55.435 ;
        RECT 186.490 55.175 186.750 55.435 ;
        RECT 183.635 54.515 183.895 54.775 ;
        RECT 186.490 54.515 186.750 54.775 ;
        RECT 183.635 53.855 183.895 54.115 ;
        RECT 186.490 53.855 186.750 54.115 ;
        RECT 183.635 53.195 183.895 53.455 ;
        RECT 186.490 53.195 186.750 53.455 ;
        RECT 183.635 52.535 183.895 52.795 ;
        RECT 186.490 52.535 186.750 52.795 ;
        RECT 183.635 51.875 183.895 52.135 ;
        RECT 186.490 51.875 186.750 52.135 ;
        RECT 183.635 51.215 183.895 51.475 ;
        RECT 186.490 51.215 186.750 51.475 ;
        RECT 183.635 50.555 183.895 50.815 ;
        RECT 186.490 50.555 186.750 50.815 ;
        RECT 182.610 22.265 182.870 22.525 ;
        RECT 182.610 21.605 182.870 21.865 ;
        RECT 182.610 20.945 182.870 21.205 ;
        RECT 183.635 18.175 183.895 18.435 ;
        RECT 186.490 18.175 186.750 18.435 ;
        RECT 183.635 17.515 183.895 17.775 ;
        RECT 186.490 17.515 186.750 17.775 ;
        RECT 183.635 16.855 183.895 17.115 ;
        RECT 186.490 16.855 186.750 17.115 ;
        RECT 183.635 16.195 183.895 16.455 ;
        RECT 186.490 16.195 186.750 16.455 ;
        RECT 183.635 15.535 183.895 15.795 ;
        RECT 186.490 15.535 186.750 15.795 ;
        RECT 183.635 14.875 183.895 15.135 ;
        RECT 186.490 14.875 186.750 15.135 ;
        RECT 183.635 14.215 183.895 14.475 ;
        RECT 186.490 14.215 186.750 14.475 ;
        RECT 183.635 13.555 183.895 13.815 ;
        RECT 186.490 13.555 186.750 13.815 ;
        RECT 183.635 12.895 183.895 13.155 ;
        RECT 186.490 12.895 186.750 13.155 ;
        RECT 183.635 12.235 183.895 12.495 ;
        RECT 186.490 12.235 186.750 12.495 ;
        RECT 183.635 11.575 183.895 11.835 ;
        RECT 186.490 11.575 186.750 11.835 ;
        RECT 183.635 10.915 183.895 11.175 ;
        RECT 186.490 10.915 186.750 11.175 ;
        RECT 183.635 10.255 183.895 10.515 ;
        RECT 186.490 10.255 186.750 10.515 ;
        RECT 183.635 9.595 183.895 9.855 ;
        RECT 186.490 9.595 186.750 9.855 ;
        RECT 183.635 8.935 183.895 9.195 ;
        RECT 186.490 8.935 186.750 9.195 ;
        RECT 188.275 55.175 188.535 55.435 ;
        RECT 191.130 55.175 191.390 55.435 ;
        RECT 188.275 54.515 188.535 54.775 ;
        RECT 191.130 54.515 191.390 54.775 ;
        RECT 188.275 53.855 188.535 54.115 ;
        RECT 191.130 53.855 191.390 54.115 ;
        RECT 188.275 53.195 188.535 53.455 ;
        RECT 191.130 53.195 191.390 53.455 ;
        RECT 188.275 52.535 188.535 52.795 ;
        RECT 191.130 52.535 191.390 52.795 ;
        RECT 188.275 51.875 188.535 52.135 ;
        RECT 191.130 51.875 191.390 52.135 ;
        RECT 188.275 51.215 188.535 51.475 ;
        RECT 191.130 51.215 191.390 51.475 ;
        RECT 188.275 50.555 188.535 50.815 ;
        RECT 191.130 50.555 191.390 50.815 ;
        RECT 187.250 24.965 187.510 25.225 ;
        RECT 187.250 24.305 187.510 24.565 ;
        RECT 187.250 23.645 187.510 23.905 ;
        RECT 188.275 18.175 188.535 18.435 ;
        RECT 191.130 18.175 191.390 18.435 ;
        RECT 188.275 17.515 188.535 17.775 ;
        RECT 191.130 17.515 191.390 17.775 ;
        RECT 188.275 16.855 188.535 17.115 ;
        RECT 191.130 16.855 191.390 17.115 ;
        RECT 188.275 16.195 188.535 16.455 ;
        RECT 191.130 16.195 191.390 16.455 ;
        RECT 188.275 15.535 188.535 15.795 ;
        RECT 191.130 15.535 191.390 15.795 ;
        RECT 188.275 14.875 188.535 15.135 ;
        RECT 191.130 14.875 191.390 15.135 ;
        RECT 188.275 14.215 188.535 14.475 ;
        RECT 191.130 14.215 191.390 14.475 ;
        RECT 188.275 13.555 188.535 13.815 ;
        RECT 191.130 13.555 191.390 13.815 ;
        RECT 188.275 12.895 188.535 13.155 ;
        RECT 191.130 12.895 191.390 13.155 ;
        RECT 188.275 12.235 188.535 12.495 ;
        RECT 191.130 12.235 191.390 12.495 ;
        RECT 188.275 11.575 188.535 11.835 ;
        RECT 191.130 11.575 191.390 11.835 ;
        RECT 188.275 10.915 188.535 11.175 ;
        RECT 191.130 10.915 191.390 11.175 ;
        RECT 188.275 10.255 188.535 10.515 ;
        RECT 191.130 10.255 191.390 10.515 ;
        RECT 188.275 9.595 188.535 9.855 ;
        RECT 191.130 9.595 191.390 9.855 ;
        RECT 188.275 8.935 188.535 9.195 ;
        RECT 191.130 8.935 191.390 9.195 ;
        RECT 192.915 55.175 193.175 55.435 ;
        RECT 192.915 54.515 193.175 54.775 ;
        RECT 192.915 53.855 193.175 54.115 ;
        RECT 192.915 53.195 193.175 53.455 ;
        RECT 192.915 52.535 193.175 52.795 ;
        RECT 192.915 51.875 193.175 52.135 ;
        RECT 192.915 51.215 193.175 51.475 ;
        RECT 192.915 50.555 193.175 50.815 ;
        RECT 191.890 45.165 192.150 45.425 ;
        RECT 191.890 44.505 192.150 44.765 ;
        RECT 191.890 43.845 192.150 44.105 ;
        RECT 192.915 18.175 193.175 18.435 ;
        RECT 192.915 17.515 193.175 17.775 ;
        RECT 192.915 16.855 193.175 17.115 ;
        RECT 192.915 16.195 193.175 16.455 ;
        RECT 192.915 15.535 193.175 15.795 ;
        RECT 192.915 14.875 193.175 15.135 ;
        RECT 192.915 14.215 193.175 14.475 ;
        RECT 192.915 13.555 193.175 13.815 ;
        RECT 192.915 12.895 193.175 13.155 ;
        RECT 192.915 12.235 193.175 12.495 ;
        RECT 192.915 11.575 193.175 11.835 ;
        RECT 192.915 10.915 193.175 11.175 ;
        RECT 192.915 10.255 193.175 10.515 ;
        RECT 192.915 9.595 193.175 9.855 ;
        RECT 192.915 8.935 193.175 9.195 ;
        RECT 4.670 8.150 4.930 8.410 ;
        RECT 4.670 7.490 4.930 7.750 ;
        RECT 4.670 6.830 4.930 7.090 ;
        RECT 0.910 4.750 1.170 5.010 ;
        RECT 2.050 4.750 2.310 5.010 ;
        RECT 3.545 4.160 3.805 4.420 ;
        RECT 22.860 8.150 23.120 8.410 ;
        RECT 22.860 7.490 23.120 7.750 ;
        RECT 22.860 6.830 23.120 7.090 ;
        RECT 8.090 4.780 8.350 5.040 ;
        RECT 8.750 4.780 9.010 5.040 ;
        RECT 9.410 4.780 9.670 5.040 ;
        RECT 14.620 4.750 14.880 5.010 ;
        RECT 15.280 4.750 15.540 5.010 ;
        RECT 15.940 4.750 16.200 5.010 ;
        RECT 17.980 4.750 18.240 5.010 ;
        RECT 18.640 4.750 18.900 5.010 ;
        RECT 19.300 4.750 19.560 5.010 ;
        RECT 4.230 3.480 4.490 3.740 ;
        RECT 4.640 2.820 4.900 3.080 ;
        RECT 7.115 3.005 7.375 3.265 ;
        RECT 9.905 2.995 10.165 3.255 ;
        RECT 3.875 2.005 4.135 2.265 ;
        RECT 0.910 0.830 1.170 1.090 ;
        RECT 2.050 0.830 2.310 1.090 ;
        RECT 7.685 2.295 7.945 2.555 ;
        RECT 11.590 2.830 12.890 3.090 ;
        RECT 15.005 2.830 15.265 3.090 ;
        RECT 12.150 1.590 12.410 1.850 ;
        RECT 16.780 1.830 17.040 2.090 ;
        RECT 20.090 3.830 20.350 4.090 ;
        RECT 21.735 4.160 21.995 4.420 ;
        RECT 42.170 8.150 42.430 8.410 ;
        RECT 42.170 7.490 42.430 7.750 ;
        RECT 42.170 6.830 42.430 7.090 ;
        RECT 26.280 4.780 26.540 5.040 ;
        RECT 26.940 4.780 27.200 5.040 ;
        RECT 27.600 4.780 27.860 5.040 ;
        RECT 32.810 4.750 33.070 5.010 ;
        RECT 33.470 4.750 33.730 5.010 ;
        RECT 34.130 4.750 34.390 5.010 ;
        RECT 36.170 4.750 36.430 5.010 ;
        RECT 36.830 4.750 37.090 5.010 ;
        RECT 37.490 4.750 37.750 5.010 ;
        RECT 39.550 4.750 39.810 5.010 ;
        RECT 22.420 3.480 22.680 3.740 ;
        RECT 18.365 2.830 18.625 3.090 ;
        RECT 22.830 2.820 23.090 3.080 ;
        RECT 25.305 3.005 25.565 3.265 ;
        RECT 28.095 2.995 28.355 3.255 ;
        RECT 22.065 2.005 22.325 2.265 ;
        RECT 7.490 0.830 7.750 1.090 ;
        RECT 8.150 0.830 8.410 1.090 ;
        RECT 8.810 0.830 9.070 1.090 ;
        RECT 14.360 0.830 14.620 1.090 ;
        RECT 15.680 0.830 15.940 1.090 ;
        RECT 17.720 0.830 17.980 1.090 ;
        RECT 19.040 0.830 19.300 1.090 ;
        RECT 25.875 2.295 26.135 2.555 ;
        RECT 29.780 2.830 31.080 3.090 ;
        RECT 33.195 2.830 33.455 3.090 ;
        RECT 30.340 1.590 30.600 1.850 ;
        RECT 34.970 1.830 35.230 2.090 ;
        RECT 38.280 3.830 38.540 4.090 ;
        RECT 41.045 4.160 41.305 4.420 ;
        RECT 57.000 8.150 57.260 8.410 ;
        RECT 57.000 7.490 57.260 7.750 ;
        RECT 57.000 6.830 57.260 7.090 ;
        RECT 45.590 4.780 45.850 5.040 ;
        RECT 46.250 4.780 46.510 5.040 ;
        RECT 46.910 4.780 47.170 5.040 ;
        RECT 52.120 4.750 52.380 5.010 ;
        RECT 52.780 4.750 53.040 5.010 ;
        RECT 53.440 4.750 53.700 5.010 ;
        RECT 41.730 3.480 41.990 3.740 ;
        RECT 36.555 2.830 36.815 3.090 ;
        RECT 42.140 2.820 42.400 3.080 ;
        RECT 44.615 3.005 44.875 3.265 ;
        RECT 47.405 2.995 47.665 3.255 ;
        RECT 41.375 2.005 41.635 2.265 ;
        RECT 25.680 0.830 25.940 1.090 ;
        RECT 26.340 0.830 26.600 1.090 ;
        RECT 27.000 0.830 27.260 1.090 ;
        RECT 32.550 0.830 32.810 1.090 ;
        RECT 33.870 0.830 34.130 1.090 ;
        RECT 35.910 0.830 36.170 1.090 ;
        RECT 37.230 0.830 37.490 1.090 ;
        RECT 39.550 0.830 39.810 1.090 ;
        RECT 45.185 2.295 45.445 2.555 ;
        RECT 49.090 2.830 50.390 3.090 ;
        RECT 55.875 4.160 56.135 4.420 ;
        RECT 60.420 4.780 60.680 5.040 ;
        RECT 61.080 4.780 61.340 5.040 ;
        RECT 61.740 4.780 62.000 5.040 ;
        RECT 66.950 4.750 67.210 5.010 ;
        RECT 67.610 4.750 67.870 5.010 ;
        RECT 68.270 4.750 68.530 5.010 ;
        RECT 70.310 4.750 70.570 5.010 ;
        RECT 70.970 4.750 71.230 5.010 ;
        RECT 71.630 4.750 71.890 5.010 ;
        RECT 73.690 4.750 73.950 5.010 ;
        RECT 74.690 4.750 74.950 5.010 ;
        RECT 75.350 4.750 75.610 5.010 ;
        RECT 76.010 4.750 76.270 5.010 ;
        RECT 76.930 4.750 77.190 5.010 ;
        RECT 77.590 4.750 77.850 5.010 ;
        RECT 78.250 4.750 78.510 5.010 ;
        RECT 79.270 4.750 79.530 5.010 ;
        RECT 79.930 4.750 80.190 5.010 ;
        RECT 80.590 4.750 80.850 5.010 ;
        RECT 82.530 4.750 82.790 5.010 ;
        RECT 83.190 4.750 83.450 5.010 ;
        RECT 83.850 4.750 84.110 5.010 ;
        RECT 84.770 4.750 85.030 5.010 ;
        RECT 85.430 4.750 85.690 5.010 ;
        RECT 86.090 4.750 86.350 5.010 ;
        RECT 87.010 4.750 87.270 5.010 ;
        RECT 87.670 4.750 87.930 5.010 ;
        RECT 88.330 4.750 88.590 5.010 ;
        RECT 89.250 4.750 89.510 5.010 ;
        RECT 89.910 4.750 90.170 5.010 ;
        RECT 90.570 4.750 90.830 5.010 ;
        RECT 91.490 4.750 91.750 5.010 ;
        RECT 92.150 4.750 92.410 5.010 ;
        RECT 92.810 4.750 93.070 5.010 ;
        RECT 93.850 4.750 94.110 5.010 ;
        RECT 94.850 4.750 95.110 5.010 ;
        RECT 95.510 4.750 95.770 5.010 ;
        RECT 96.170 4.750 96.430 5.010 ;
        RECT 97.090 4.750 97.350 5.010 ;
        RECT 97.750 4.750 98.010 5.010 ;
        RECT 98.410 4.750 98.670 5.010 ;
        RECT 99.330 4.750 99.590 5.010 ;
        RECT 99.990 4.750 100.250 5.010 ;
        RECT 100.650 4.750 100.910 5.010 ;
        RECT 101.670 4.750 101.930 5.010 ;
        RECT 102.330 4.750 102.590 5.010 ;
        RECT 102.990 4.750 103.250 5.010 ;
        RECT 104.930 4.750 105.190 5.010 ;
        RECT 105.590 4.750 105.850 5.010 ;
        RECT 106.250 4.750 106.510 5.010 ;
        RECT 107.170 4.750 107.430 5.010 ;
        RECT 107.830 4.750 108.090 5.010 ;
        RECT 108.490 4.750 108.750 5.010 ;
        RECT 109.410 4.750 109.670 5.010 ;
        RECT 110.070 4.750 110.330 5.010 ;
        RECT 110.730 4.750 110.990 5.010 ;
        RECT 111.650 4.750 111.910 5.010 ;
        RECT 112.310 4.750 112.570 5.010 ;
        RECT 112.970 4.750 113.230 5.010 ;
        RECT 114.010 4.750 114.270 5.010 ;
        RECT 115.010 4.750 115.270 5.010 ;
        RECT 115.670 4.750 115.930 5.010 ;
        RECT 116.330 4.750 116.590 5.010 ;
        RECT 117.250 4.750 117.510 5.010 ;
        RECT 117.910 4.750 118.170 5.010 ;
        RECT 118.570 4.750 118.830 5.010 ;
        RECT 119.490 4.750 119.750 5.010 ;
        RECT 120.150 4.750 120.410 5.010 ;
        RECT 120.810 4.750 121.070 5.010 ;
        RECT 121.830 4.750 122.090 5.010 ;
        RECT 122.490 4.750 122.750 5.010 ;
        RECT 123.150 4.750 123.410 5.010 ;
        RECT 125.090 4.750 125.350 5.010 ;
        RECT 125.750 4.750 126.010 5.010 ;
        RECT 126.410 4.750 126.670 5.010 ;
        RECT 127.330 4.750 127.590 5.010 ;
        RECT 127.990 4.750 128.250 5.010 ;
        RECT 128.650 4.750 128.910 5.010 ;
        RECT 129.570 4.750 129.830 5.010 ;
        RECT 130.230 4.750 130.490 5.010 ;
        RECT 130.890 4.750 131.150 5.010 ;
        RECT 131.810 4.750 132.070 5.010 ;
        RECT 132.470 4.750 132.730 5.010 ;
        RECT 133.130 4.750 133.390 5.010 ;
        RECT 134.170 4.750 134.430 5.010 ;
        RECT 135.170 4.750 135.430 5.010 ;
        RECT 135.830 4.750 136.090 5.010 ;
        RECT 136.490 4.750 136.750 5.010 ;
        RECT 137.410 4.750 137.670 5.010 ;
        RECT 138.070 4.750 138.330 5.010 ;
        RECT 138.730 4.750 138.990 5.010 ;
        RECT 139.650 4.750 139.910 5.010 ;
        RECT 140.310 4.750 140.570 5.010 ;
        RECT 140.970 4.750 141.230 5.010 ;
        RECT 141.890 4.750 142.150 5.010 ;
        RECT 142.550 4.750 142.810 5.010 ;
        RECT 143.210 4.750 143.470 5.010 ;
        RECT 144.230 4.750 144.490 5.010 ;
        RECT 144.890 4.750 145.150 5.010 ;
        RECT 145.550 4.750 145.810 5.010 ;
        RECT 147.490 4.750 147.750 5.010 ;
        RECT 148.150 4.750 148.410 5.010 ;
        RECT 148.810 4.750 149.070 5.010 ;
        RECT 149.730 4.750 149.990 5.010 ;
        RECT 150.390 4.750 150.650 5.010 ;
        RECT 151.050 4.750 151.310 5.010 ;
        RECT 151.970 4.750 152.230 5.010 ;
        RECT 152.630 4.750 152.890 5.010 ;
        RECT 153.290 4.750 153.550 5.010 ;
        RECT 154.330 4.750 154.590 5.010 ;
        RECT 155.330 4.750 155.590 5.010 ;
        RECT 155.990 4.750 156.250 5.010 ;
        RECT 156.650 4.750 156.910 5.010 ;
        RECT 157.570 4.750 157.830 5.010 ;
        RECT 158.230 4.750 158.490 5.010 ;
        RECT 158.890 4.750 159.150 5.010 ;
        RECT 159.810 4.750 160.070 5.010 ;
        RECT 160.470 4.750 160.730 5.010 ;
        RECT 161.130 4.750 161.390 5.010 ;
        RECT 162.050 4.750 162.310 5.010 ;
        RECT 162.710 4.750 162.970 5.010 ;
        RECT 163.370 4.750 163.630 5.010 ;
        RECT 164.290 4.750 164.550 5.010 ;
        RECT 164.950 4.750 165.210 5.010 ;
        RECT 165.610 4.750 165.870 5.010 ;
        RECT 166.630 4.750 166.890 5.010 ;
        RECT 167.290 4.750 167.550 5.010 ;
        RECT 167.950 4.750 168.210 5.010 ;
        RECT 169.890 4.750 170.150 5.010 ;
        RECT 170.550 4.750 170.810 5.010 ;
        RECT 171.210 4.750 171.470 5.010 ;
        RECT 172.130 4.750 172.390 5.010 ;
        RECT 172.790 4.750 173.050 5.010 ;
        RECT 173.450 4.750 173.710 5.010 ;
        RECT 174.470 4.750 174.730 5.010 ;
        RECT 56.560 3.480 56.820 3.740 ;
        RECT 52.505 2.830 52.765 3.090 ;
        RECT 56.970 2.820 57.230 3.080 ;
        RECT 59.445 3.005 59.705 3.265 ;
        RECT 62.235 2.995 62.495 3.255 ;
        RECT 49.650 1.590 49.910 1.850 ;
        RECT 54.280 1.830 54.540 2.090 ;
        RECT 56.205 2.005 56.465 2.265 ;
        RECT 44.990 0.830 45.250 1.090 ;
        RECT 45.650 0.830 45.910 1.090 ;
        RECT 46.310 0.830 46.570 1.090 ;
        RECT 51.860 0.830 52.120 1.090 ;
        RECT 53.180 0.830 53.440 1.090 ;
        RECT 60.015 2.295 60.275 2.555 ;
        RECT 63.920 2.830 65.220 3.090 ;
        RECT 67.335 2.830 67.595 3.090 ;
        RECT 64.480 1.590 64.740 1.850 ;
        RECT 69.110 1.830 69.370 2.090 ;
        RECT 72.420 3.830 72.680 4.090 ;
        RECT 70.695 2.830 70.955 3.090 ;
        RECT 81.380 3.830 81.640 4.090 ;
        RECT 79.655 2.830 79.915 3.090 ;
        RECT 103.780 3.830 104.040 4.090 ;
        RECT 102.055 2.830 102.315 3.090 ;
        RECT 123.940 3.830 124.200 4.090 ;
        RECT 122.215 2.830 122.475 3.090 ;
        RECT 146.340 3.830 146.600 4.090 ;
        RECT 144.615 2.830 144.875 3.090 ;
        RECT 168.740 3.830 169.000 4.090 ;
        RECT 167.015 2.830 167.275 3.090 ;
        RECT 59.820 0.830 60.080 1.090 ;
        RECT 60.480 0.830 60.740 1.090 ;
        RECT 61.140 0.830 61.400 1.090 ;
        RECT 66.690 0.830 66.950 1.090 ;
        RECT 68.010 0.830 68.270 1.090 ;
        RECT 70.050 0.830 70.310 1.090 ;
        RECT 71.370 0.830 71.630 1.090 ;
        RECT 73.690 0.830 73.950 1.090 ;
        RECT 74.690 0.830 74.950 1.090 ;
        RECT 75.350 0.830 75.610 1.090 ;
        RECT 76.010 0.830 76.270 1.090 ;
        RECT 76.930 0.830 77.190 1.090 ;
        RECT 77.590 0.830 77.850 1.090 ;
        RECT 78.250 0.830 78.510 1.090 ;
        RECT 79.010 0.830 79.270 1.090 ;
        RECT 80.330 0.830 80.590 1.090 ;
        RECT 82.530 0.830 82.790 1.090 ;
        RECT 83.190 0.830 83.450 1.090 ;
        RECT 83.850 0.830 84.110 1.090 ;
        RECT 84.770 0.830 85.030 1.090 ;
        RECT 85.430 0.830 85.690 1.090 ;
        RECT 86.090 0.830 86.350 1.090 ;
        RECT 87.010 0.830 87.270 1.090 ;
        RECT 87.670 0.830 87.930 1.090 ;
        RECT 88.330 0.830 88.590 1.090 ;
        RECT 89.250 0.830 89.510 1.090 ;
        RECT 89.910 0.830 90.170 1.090 ;
        RECT 90.570 0.830 90.830 1.090 ;
        RECT 91.490 0.830 91.750 1.090 ;
        RECT 92.150 0.830 92.410 1.090 ;
        RECT 92.810 0.830 93.070 1.090 ;
        RECT 93.850 0.830 94.110 1.090 ;
        RECT 94.850 0.830 95.110 1.090 ;
        RECT 95.510 0.830 95.770 1.090 ;
        RECT 96.170 0.830 96.430 1.090 ;
        RECT 97.090 0.830 97.350 1.090 ;
        RECT 97.750 0.830 98.010 1.090 ;
        RECT 98.410 0.830 98.670 1.090 ;
        RECT 99.330 0.830 99.590 1.090 ;
        RECT 99.990 0.830 100.250 1.090 ;
        RECT 100.650 0.830 100.910 1.090 ;
        RECT 101.410 0.830 101.670 1.090 ;
        RECT 102.730 0.830 102.990 1.090 ;
        RECT 104.930 0.830 105.190 1.090 ;
        RECT 105.590 0.830 105.850 1.090 ;
        RECT 106.250 0.830 106.510 1.090 ;
        RECT 107.170 0.830 107.430 1.090 ;
        RECT 107.830 0.830 108.090 1.090 ;
        RECT 108.490 0.830 108.750 1.090 ;
        RECT 109.410 0.830 109.670 1.090 ;
        RECT 110.070 0.830 110.330 1.090 ;
        RECT 110.730 0.830 110.990 1.090 ;
        RECT 111.650 0.830 111.910 1.090 ;
        RECT 112.310 0.830 112.570 1.090 ;
        RECT 112.970 0.830 113.230 1.090 ;
        RECT 114.010 0.830 114.270 1.090 ;
        RECT 115.010 0.830 115.270 1.090 ;
        RECT 115.670 0.830 115.930 1.090 ;
        RECT 116.330 0.830 116.590 1.090 ;
        RECT 117.250 0.830 117.510 1.090 ;
        RECT 117.910 0.830 118.170 1.090 ;
        RECT 118.570 0.830 118.830 1.090 ;
        RECT 119.490 0.830 119.750 1.090 ;
        RECT 120.150 0.830 120.410 1.090 ;
        RECT 120.810 0.830 121.070 1.090 ;
        RECT 121.570 0.830 121.830 1.090 ;
        RECT 122.890 0.830 123.150 1.090 ;
        RECT 125.090 0.830 125.350 1.090 ;
        RECT 125.750 0.830 126.010 1.090 ;
        RECT 126.410 0.830 126.670 1.090 ;
        RECT 127.330 0.830 127.590 1.090 ;
        RECT 127.990 0.830 128.250 1.090 ;
        RECT 128.650 0.830 128.910 1.090 ;
        RECT 129.570 0.830 129.830 1.090 ;
        RECT 130.230 0.830 130.490 1.090 ;
        RECT 130.890 0.830 131.150 1.090 ;
        RECT 131.810 0.830 132.070 1.090 ;
        RECT 132.470 0.830 132.730 1.090 ;
        RECT 133.130 0.830 133.390 1.090 ;
        RECT 134.170 0.830 134.430 1.090 ;
        RECT 135.170 0.830 135.430 1.090 ;
        RECT 135.830 0.830 136.090 1.090 ;
        RECT 136.490 0.830 136.750 1.090 ;
        RECT 137.410 0.830 137.670 1.090 ;
        RECT 138.070 0.830 138.330 1.090 ;
        RECT 138.730 0.830 138.990 1.090 ;
        RECT 139.650 0.830 139.910 1.090 ;
        RECT 140.310 0.830 140.570 1.090 ;
        RECT 140.970 0.830 141.230 1.090 ;
        RECT 141.890 0.830 142.150 1.090 ;
        RECT 142.550 0.830 142.810 1.090 ;
        RECT 143.210 0.830 143.470 1.090 ;
        RECT 143.970 0.830 144.230 1.090 ;
        RECT 145.290 0.830 145.550 1.090 ;
        RECT 147.490 0.830 147.750 1.090 ;
        RECT 148.150 0.830 148.410 1.090 ;
        RECT 148.810 0.830 149.070 1.090 ;
        RECT 149.730 0.830 149.990 1.090 ;
        RECT 150.390 0.830 150.650 1.090 ;
        RECT 151.050 0.830 151.310 1.090 ;
        RECT 151.970 0.830 152.230 1.090 ;
        RECT 152.630 0.830 152.890 1.090 ;
        RECT 153.290 0.830 153.550 1.090 ;
        RECT 154.330 0.830 154.590 1.090 ;
        RECT 155.330 0.830 155.590 1.090 ;
        RECT 155.990 0.830 156.250 1.090 ;
        RECT 156.650 0.830 156.910 1.090 ;
        RECT 157.570 0.830 157.830 1.090 ;
        RECT 158.230 0.830 158.490 1.090 ;
        RECT 158.890 0.830 159.150 1.090 ;
        RECT 159.810 0.830 160.070 1.090 ;
        RECT 160.470 0.830 160.730 1.090 ;
        RECT 161.130 0.830 161.390 1.090 ;
        RECT 162.050 0.830 162.310 1.090 ;
        RECT 162.710 0.830 162.970 1.090 ;
        RECT 163.370 0.830 163.630 1.090 ;
        RECT 164.290 0.830 164.550 1.090 ;
        RECT 164.950 0.830 165.210 1.090 ;
        RECT 165.610 0.830 165.870 1.090 ;
        RECT 166.370 0.830 166.630 1.090 ;
        RECT 167.690 0.830 167.950 1.090 ;
        RECT 169.890 0.830 170.150 1.090 ;
        RECT 170.550 0.830 170.810 1.090 ;
        RECT 171.210 0.830 171.470 1.090 ;
        RECT 172.130 0.830 172.390 1.090 ;
        RECT 172.790 0.830 173.050 1.090 ;
        RECT 173.450 0.830 173.710 1.090 ;
        RECT 174.470 0.830 174.730 1.090 ;
      LAYER Metal2 ;
        RECT 1.975 59.890 20.510 60.305 ;
        RECT 23.970 59.890 42.505 60.305 ;
        RECT 45.965 59.890 64.500 60.305 ;
        RECT 67.960 59.890 86.495 60.305 ;
        RECT 89.955 59.890 108.490 60.305 ;
        RECT 111.950 59.890 130.485 60.305 ;
        RECT 133.945 59.890 152.480 60.305 ;
        RECT 155.940 59.890 174.475 60.305 ;
        RECT 0.765 58.745 1.145 59.125 ;
        RECT 0.765 58.085 1.145 58.465 ;
        RECT 0.765 57.425 1.145 57.805 ;
        RECT 0.765 56.765 1.145 57.145 ;
        RECT 0.765 56.105 1.145 56.485 ;
        RECT 0.765 55.445 1.145 55.825 ;
        RECT 0.765 54.785 1.145 55.165 ;
        RECT 0.765 54.125 1.145 54.505 ;
        RECT 0.765 53.465 1.145 53.845 ;
        RECT 0.765 52.805 1.145 53.185 ;
        RECT 0.765 52.145 1.145 52.525 ;
        RECT 0.765 51.485 1.145 51.865 ;
        RECT 0.765 50.825 1.145 51.205 ;
        RECT 0.765 50.165 1.145 50.545 ;
        RECT 5.250 47.805 5.630 48.185 ;
        RECT 5.910 47.805 6.290 48.185 ;
        RECT 6.570 47.805 6.950 48.185 ;
        RECT 5.250 47.145 5.630 47.525 ;
        RECT 5.910 47.145 6.290 47.525 ;
        RECT 6.570 47.145 6.950 47.525 ;
        RECT 5.250 46.485 5.630 46.865 ;
        RECT 5.910 46.485 6.290 46.865 ;
        RECT 6.570 46.485 6.950 46.865 ;
        RECT 5.250 22.205 5.630 22.585 ;
        RECT 5.910 22.205 6.290 22.585 ;
        RECT 6.570 22.205 6.950 22.585 ;
        RECT 5.250 21.545 5.630 21.925 ;
        RECT 5.910 21.545 6.290 21.925 ;
        RECT 6.570 21.545 6.950 21.925 ;
        RECT 5.250 20.885 5.630 21.265 ;
        RECT 5.910 20.885 6.290 21.265 ;
        RECT 6.570 20.885 6.950 21.265 ;
        RECT 9.000 9.150 9.525 59.890 ;
        RECT 11.055 58.745 11.435 59.125 ;
        RECT 11.055 58.085 11.435 58.465 ;
        RECT 11.055 57.425 11.435 57.805 ;
        RECT 11.055 56.765 11.435 57.145 ;
        RECT 11.055 56.105 11.435 56.485 ;
        RECT 11.055 55.445 11.435 55.825 ;
        RECT 11.055 54.785 11.435 55.165 ;
        RECT 11.055 54.125 11.435 54.505 ;
        RECT 11.055 53.465 11.435 53.845 ;
        RECT 11.055 52.805 11.435 53.185 ;
        RECT 11.055 52.145 11.435 52.525 ;
        RECT 11.055 51.485 11.435 51.865 ;
        RECT 11.055 50.825 11.435 51.205 ;
        RECT 11.055 50.165 11.435 50.545 ;
        RECT 12.440 9.150 12.965 59.890 ;
        RECT 21.340 58.745 21.720 59.125 ;
        RECT 22.760 58.745 23.140 59.125 ;
        RECT 21.340 58.085 21.720 58.465 ;
        RECT 22.760 58.085 23.140 58.465 ;
        RECT 21.340 57.425 21.720 57.805 ;
        RECT 22.760 57.425 23.140 57.805 ;
        RECT 21.340 56.765 21.720 57.145 ;
        RECT 22.760 56.765 23.140 57.145 ;
        RECT 21.340 56.105 21.720 56.485 ;
        RECT 22.760 56.105 23.140 56.485 ;
        RECT 21.340 55.445 21.720 55.825 ;
        RECT 22.760 55.445 23.140 55.825 ;
        RECT 21.340 54.785 21.720 55.165 ;
        RECT 22.760 54.785 23.140 55.165 ;
        RECT 21.340 54.125 21.720 54.505 ;
        RECT 22.760 54.125 23.140 54.505 ;
        RECT 21.340 53.465 21.720 53.845 ;
        RECT 22.760 53.465 23.140 53.845 ;
        RECT 21.340 52.805 21.720 53.185 ;
        RECT 22.760 52.805 23.140 53.185 ;
        RECT 21.340 52.145 21.720 52.525 ;
        RECT 22.760 52.145 23.140 52.525 ;
        RECT 21.340 51.485 21.720 51.865 ;
        RECT 22.760 51.485 23.140 51.865 ;
        RECT 21.340 50.825 21.720 51.205 ;
        RECT 22.760 50.825 23.140 51.205 ;
        RECT 21.340 50.165 21.720 50.545 ;
        RECT 22.760 50.165 23.140 50.545 ;
        RECT 27.245 47.805 27.625 48.185 ;
        RECT 27.905 47.805 28.285 48.185 ;
        RECT 28.565 47.805 28.945 48.185 ;
        RECT 27.245 47.145 27.625 47.525 ;
        RECT 27.905 47.145 28.285 47.525 ;
        RECT 28.565 47.145 28.945 47.525 ;
        RECT 27.245 46.485 27.625 46.865 ;
        RECT 27.905 46.485 28.285 46.865 ;
        RECT 28.565 46.485 28.945 46.865 ;
        RECT 15.550 45.105 15.930 45.485 ;
        RECT 16.210 45.105 16.590 45.485 ;
        RECT 16.870 45.105 17.250 45.485 ;
        RECT 15.550 44.445 15.930 44.825 ;
        RECT 16.210 44.445 16.590 44.825 ;
        RECT 16.870 44.445 17.250 44.825 ;
        RECT 15.550 43.785 15.930 44.165 ;
        RECT 16.210 43.785 16.590 44.165 ;
        RECT 16.870 43.785 17.250 44.165 ;
        RECT 15.550 24.905 15.930 25.285 ;
        RECT 16.210 24.905 16.590 25.285 ;
        RECT 16.870 24.905 17.250 25.285 ;
        RECT 15.550 24.245 15.930 24.625 ;
        RECT 16.210 24.245 16.590 24.625 ;
        RECT 16.870 24.245 17.250 24.625 ;
        RECT 15.550 23.585 15.930 23.965 ;
        RECT 16.210 23.585 16.590 23.965 ;
        RECT 16.870 23.585 17.250 23.965 ;
        RECT 27.245 22.205 27.625 22.585 ;
        RECT 27.905 22.205 28.285 22.585 ;
        RECT 28.565 22.205 28.945 22.585 ;
        RECT 27.245 21.545 27.625 21.925 ;
        RECT 27.905 21.545 28.285 21.925 ;
        RECT 28.565 21.545 28.945 21.925 ;
        RECT 27.245 20.885 27.625 21.265 ;
        RECT 27.905 20.885 28.285 21.265 ;
        RECT 28.565 20.885 28.945 21.265 ;
        RECT 9.000 9.100 12.965 9.150 ;
        RECT 30.995 9.150 31.520 59.890 ;
        RECT 33.050 58.745 33.430 59.125 ;
        RECT 33.050 58.085 33.430 58.465 ;
        RECT 33.050 57.425 33.430 57.805 ;
        RECT 33.050 56.765 33.430 57.145 ;
        RECT 33.050 56.105 33.430 56.485 ;
        RECT 33.050 55.445 33.430 55.825 ;
        RECT 33.050 54.785 33.430 55.165 ;
        RECT 33.050 54.125 33.430 54.505 ;
        RECT 33.050 53.465 33.430 53.845 ;
        RECT 33.050 52.805 33.430 53.185 ;
        RECT 33.050 52.145 33.430 52.525 ;
        RECT 33.050 51.485 33.430 51.865 ;
        RECT 33.050 50.825 33.430 51.205 ;
        RECT 33.050 50.165 33.430 50.545 ;
        RECT 34.435 9.150 34.960 59.890 ;
        RECT 43.335 58.745 43.715 59.125 ;
        RECT 44.755 58.745 45.135 59.125 ;
        RECT 43.335 58.085 43.715 58.465 ;
        RECT 44.755 58.085 45.135 58.465 ;
        RECT 43.335 57.425 43.715 57.805 ;
        RECT 44.755 57.425 45.135 57.805 ;
        RECT 43.335 56.765 43.715 57.145 ;
        RECT 44.755 56.765 45.135 57.145 ;
        RECT 43.335 56.105 43.715 56.485 ;
        RECT 44.755 56.105 45.135 56.485 ;
        RECT 43.335 55.445 43.715 55.825 ;
        RECT 44.755 55.445 45.135 55.825 ;
        RECT 43.335 54.785 43.715 55.165 ;
        RECT 44.755 54.785 45.135 55.165 ;
        RECT 43.335 54.125 43.715 54.505 ;
        RECT 44.755 54.125 45.135 54.505 ;
        RECT 43.335 53.465 43.715 53.845 ;
        RECT 44.755 53.465 45.135 53.845 ;
        RECT 43.335 52.805 43.715 53.185 ;
        RECT 44.755 52.805 45.135 53.185 ;
        RECT 43.335 52.145 43.715 52.525 ;
        RECT 44.755 52.145 45.135 52.525 ;
        RECT 43.335 51.485 43.715 51.865 ;
        RECT 44.755 51.485 45.135 51.865 ;
        RECT 43.335 50.825 43.715 51.205 ;
        RECT 44.755 50.825 45.135 51.205 ;
        RECT 43.335 50.165 43.715 50.545 ;
        RECT 44.755 50.165 45.135 50.545 ;
        RECT 49.240 47.805 49.620 48.185 ;
        RECT 49.900 47.805 50.280 48.185 ;
        RECT 50.560 47.805 50.940 48.185 ;
        RECT 49.240 47.145 49.620 47.525 ;
        RECT 49.900 47.145 50.280 47.525 ;
        RECT 50.560 47.145 50.940 47.525 ;
        RECT 49.240 46.485 49.620 46.865 ;
        RECT 49.900 46.485 50.280 46.865 ;
        RECT 50.560 46.485 50.940 46.865 ;
        RECT 37.545 45.105 37.925 45.485 ;
        RECT 38.205 45.105 38.585 45.485 ;
        RECT 38.865 45.105 39.245 45.485 ;
        RECT 37.545 44.445 37.925 44.825 ;
        RECT 38.205 44.445 38.585 44.825 ;
        RECT 38.865 44.445 39.245 44.825 ;
        RECT 37.545 43.785 37.925 44.165 ;
        RECT 38.205 43.785 38.585 44.165 ;
        RECT 38.865 43.785 39.245 44.165 ;
        RECT 37.545 24.905 37.925 25.285 ;
        RECT 38.205 24.905 38.585 25.285 ;
        RECT 38.865 24.905 39.245 25.285 ;
        RECT 37.545 24.245 37.925 24.625 ;
        RECT 38.205 24.245 38.585 24.625 ;
        RECT 38.865 24.245 39.245 24.625 ;
        RECT 37.545 23.585 37.925 23.965 ;
        RECT 38.205 23.585 38.585 23.965 ;
        RECT 38.865 23.585 39.245 23.965 ;
        RECT 49.240 22.205 49.620 22.585 ;
        RECT 49.900 22.205 50.280 22.585 ;
        RECT 50.560 22.205 50.940 22.585 ;
        RECT 49.240 21.545 49.620 21.925 ;
        RECT 49.900 21.545 50.280 21.925 ;
        RECT 50.560 21.545 50.940 21.925 ;
        RECT 49.240 20.885 49.620 21.265 ;
        RECT 49.900 20.885 50.280 21.265 ;
        RECT 50.560 20.885 50.940 21.265 ;
        RECT 30.995 9.100 34.960 9.150 ;
        RECT 52.990 9.150 53.515 59.890 ;
        RECT 55.045 58.745 55.425 59.125 ;
        RECT 55.045 58.085 55.425 58.465 ;
        RECT 55.045 57.425 55.425 57.805 ;
        RECT 55.045 56.765 55.425 57.145 ;
        RECT 55.045 56.105 55.425 56.485 ;
        RECT 55.045 55.445 55.425 55.825 ;
        RECT 55.045 54.785 55.425 55.165 ;
        RECT 55.045 54.125 55.425 54.505 ;
        RECT 55.045 53.465 55.425 53.845 ;
        RECT 55.045 52.805 55.425 53.185 ;
        RECT 55.045 52.145 55.425 52.525 ;
        RECT 55.045 51.485 55.425 51.865 ;
        RECT 55.045 50.825 55.425 51.205 ;
        RECT 55.045 50.165 55.425 50.545 ;
        RECT 56.430 9.150 56.955 59.890 ;
        RECT 65.330 58.745 65.710 59.125 ;
        RECT 66.750 58.745 67.130 59.125 ;
        RECT 65.330 58.085 65.710 58.465 ;
        RECT 66.750 58.085 67.130 58.465 ;
        RECT 65.330 57.425 65.710 57.805 ;
        RECT 66.750 57.425 67.130 57.805 ;
        RECT 65.330 56.765 65.710 57.145 ;
        RECT 66.750 56.765 67.130 57.145 ;
        RECT 65.330 56.105 65.710 56.485 ;
        RECT 66.750 56.105 67.130 56.485 ;
        RECT 65.330 55.445 65.710 55.825 ;
        RECT 66.750 55.445 67.130 55.825 ;
        RECT 65.330 54.785 65.710 55.165 ;
        RECT 66.750 54.785 67.130 55.165 ;
        RECT 65.330 54.125 65.710 54.505 ;
        RECT 66.750 54.125 67.130 54.505 ;
        RECT 65.330 53.465 65.710 53.845 ;
        RECT 66.750 53.465 67.130 53.845 ;
        RECT 65.330 52.805 65.710 53.185 ;
        RECT 66.750 52.805 67.130 53.185 ;
        RECT 65.330 52.145 65.710 52.525 ;
        RECT 66.750 52.145 67.130 52.525 ;
        RECT 65.330 51.485 65.710 51.865 ;
        RECT 66.750 51.485 67.130 51.865 ;
        RECT 65.330 50.825 65.710 51.205 ;
        RECT 66.750 50.825 67.130 51.205 ;
        RECT 65.330 50.165 65.710 50.545 ;
        RECT 66.750 50.165 67.130 50.545 ;
        RECT 71.235 47.805 71.615 48.185 ;
        RECT 71.895 47.805 72.275 48.185 ;
        RECT 72.555 47.805 72.935 48.185 ;
        RECT 71.235 47.145 71.615 47.525 ;
        RECT 71.895 47.145 72.275 47.525 ;
        RECT 72.555 47.145 72.935 47.525 ;
        RECT 71.235 46.485 71.615 46.865 ;
        RECT 71.895 46.485 72.275 46.865 ;
        RECT 72.555 46.485 72.935 46.865 ;
        RECT 59.540 45.105 59.920 45.485 ;
        RECT 60.200 45.105 60.580 45.485 ;
        RECT 60.860 45.105 61.240 45.485 ;
        RECT 59.540 44.445 59.920 44.825 ;
        RECT 60.200 44.445 60.580 44.825 ;
        RECT 60.860 44.445 61.240 44.825 ;
        RECT 59.540 43.785 59.920 44.165 ;
        RECT 60.200 43.785 60.580 44.165 ;
        RECT 60.860 43.785 61.240 44.165 ;
        RECT 59.540 24.905 59.920 25.285 ;
        RECT 60.200 24.905 60.580 25.285 ;
        RECT 60.860 24.905 61.240 25.285 ;
        RECT 59.540 24.245 59.920 24.625 ;
        RECT 60.200 24.245 60.580 24.625 ;
        RECT 60.860 24.245 61.240 24.625 ;
        RECT 59.540 23.585 59.920 23.965 ;
        RECT 60.200 23.585 60.580 23.965 ;
        RECT 60.860 23.585 61.240 23.965 ;
        RECT 71.235 22.205 71.615 22.585 ;
        RECT 71.895 22.205 72.275 22.585 ;
        RECT 72.555 22.205 72.935 22.585 ;
        RECT 71.235 21.545 71.615 21.925 ;
        RECT 71.895 21.545 72.275 21.925 ;
        RECT 72.555 21.545 72.935 21.925 ;
        RECT 71.235 20.885 71.615 21.265 ;
        RECT 71.895 20.885 72.275 21.265 ;
        RECT 72.555 20.885 72.935 21.265 ;
        RECT 52.990 9.100 56.955 9.150 ;
        RECT 74.985 9.150 75.510 59.890 ;
        RECT 77.040 58.745 77.420 59.125 ;
        RECT 77.040 58.085 77.420 58.465 ;
        RECT 77.040 57.425 77.420 57.805 ;
        RECT 77.040 56.765 77.420 57.145 ;
        RECT 77.040 56.105 77.420 56.485 ;
        RECT 77.040 55.445 77.420 55.825 ;
        RECT 77.040 54.785 77.420 55.165 ;
        RECT 77.040 54.125 77.420 54.505 ;
        RECT 77.040 53.465 77.420 53.845 ;
        RECT 77.040 52.805 77.420 53.185 ;
        RECT 77.040 52.145 77.420 52.525 ;
        RECT 77.040 51.485 77.420 51.865 ;
        RECT 77.040 50.825 77.420 51.205 ;
        RECT 77.040 50.165 77.420 50.545 ;
        RECT 78.425 9.150 78.950 59.890 ;
        RECT 87.325 58.745 87.705 59.125 ;
        RECT 88.745 58.745 89.125 59.125 ;
        RECT 87.325 58.085 87.705 58.465 ;
        RECT 88.745 58.085 89.125 58.465 ;
        RECT 87.325 57.425 87.705 57.805 ;
        RECT 88.745 57.425 89.125 57.805 ;
        RECT 87.325 56.765 87.705 57.145 ;
        RECT 88.745 56.765 89.125 57.145 ;
        RECT 87.325 56.105 87.705 56.485 ;
        RECT 88.745 56.105 89.125 56.485 ;
        RECT 87.325 55.445 87.705 55.825 ;
        RECT 88.745 55.445 89.125 55.825 ;
        RECT 87.325 54.785 87.705 55.165 ;
        RECT 88.745 54.785 89.125 55.165 ;
        RECT 87.325 54.125 87.705 54.505 ;
        RECT 88.745 54.125 89.125 54.505 ;
        RECT 87.325 53.465 87.705 53.845 ;
        RECT 88.745 53.465 89.125 53.845 ;
        RECT 87.325 52.805 87.705 53.185 ;
        RECT 88.745 52.805 89.125 53.185 ;
        RECT 87.325 52.145 87.705 52.525 ;
        RECT 88.745 52.145 89.125 52.525 ;
        RECT 87.325 51.485 87.705 51.865 ;
        RECT 88.745 51.485 89.125 51.865 ;
        RECT 87.325 50.825 87.705 51.205 ;
        RECT 88.745 50.825 89.125 51.205 ;
        RECT 87.325 50.165 87.705 50.545 ;
        RECT 88.745 50.165 89.125 50.545 ;
        RECT 93.230 47.805 93.610 48.185 ;
        RECT 93.890 47.805 94.270 48.185 ;
        RECT 94.550 47.805 94.930 48.185 ;
        RECT 93.230 47.145 93.610 47.525 ;
        RECT 93.890 47.145 94.270 47.525 ;
        RECT 94.550 47.145 94.930 47.525 ;
        RECT 93.230 46.485 93.610 46.865 ;
        RECT 93.890 46.485 94.270 46.865 ;
        RECT 94.550 46.485 94.930 46.865 ;
        RECT 81.535 45.105 81.915 45.485 ;
        RECT 82.195 45.105 82.575 45.485 ;
        RECT 82.855 45.105 83.235 45.485 ;
        RECT 81.535 44.445 81.915 44.825 ;
        RECT 82.195 44.445 82.575 44.825 ;
        RECT 82.855 44.445 83.235 44.825 ;
        RECT 81.535 43.785 81.915 44.165 ;
        RECT 82.195 43.785 82.575 44.165 ;
        RECT 82.855 43.785 83.235 44.165 ;
        RECT 81.535 24.905 81.915 25.285 ;
        RECT 82.195 24.905 82.575 25.285 ;
        RECT 82.855 24.905 83.235 25.285 ;
        RECT 81.535 24.245 81.915 24.625 ;
        RECT 82.195 24.245 82.575 24.625 ;
        RECT 82.855 24.245 83.235 24.625 ;
        RECT 81.535 23.585 81.915 23.965 ;
        RECT 82.195 23.585 82.575 23.965 ;
        RECT 82.855 23.585 83.235 23.965 ;
        RECT 93.230 22.205 93.610 22.585 ;
        RECT 93.890 22.205 94.270 22.585 ;
        RECT 94.550 22.205 94.930 22.585 ;
        RECT 93.230 21.545 93.610 21.925 ;
        RECT 93.890 21.545 94.270 21.925 ;
        RECT 94.550 21.545 94.930 21.925 ;
        RECT 93.230 20.885 93.610 21.265 ;
        RECT 93.890 20.885 94.270 21.265 ;
        RECT 94.550 20.885 94.930 21.265 ;
        RECT 74.985 9.100 78.950 9.150 ;
        RECT 96.980 9.150 97.505 59.890 ;
        RECT 99.035 58.745 99.415 59.125 ;
        RECT 99.035 58.085 99.415 58.465 ;
        RECT 99.035 57.425 99.415 57.805 ;
        RECT 99.035 56.765 99.415 57.145 ;
        RECT 99.035 56.105 99.415 56.485 ;
        RECT 99.035 55.445 99.415 55.825 ;
        RECT 99.035 54.785 99.415 55.165 ;
        RECT 99.035 54.125 99.415 54.505 ;
        RECT 99.035 53.465 99.415 53.845 ;
        RECT 99.035 52.805 99.415 53.185 ;
        RECT 99.035 52.145 99.415 52.525 ;
        RECT 99.035 51.485 99.415 51.865 ;
        RECT 99.035 50.825 99.415 51.205 ;
        RECT 99.035 50.165 99.415 50.545 ;
        RECT 100.420 9.150 100.945 59.890 ;
        RECT 109.320 58.745 109.700 59.125 ;
        RECT 110.740 58.745 111.120 59.125 ;
        RECT 109.320 58.085 109.700 58.465 ;
        RECT 110.740 58.085 111.120 58.465 ;
        RECT 109.320 57.425 109.700 57.805 ;
        RECT 110.740 57.425 111.120 57.805 ;
        RECT 109.320 56.765 109.700 57.145 ;
        RECT 110.740 56.765 111.120 57.145 ;
        RECT 109.320 56.105 109.700 56.485 ;
        RECT 110.740 56.105 111.120 56.485 ;
        RECT 109.320 55.445 109.700 55.825 ;
        RECT 110.740 55.445 111.120 55.825 ;
        RECT 109.320 54.785 109.700 55.165 ;
        RECT 110.740 54.785 111.120 55.165 ;
        RECT 109.320 54.125 109.700 54.505 ;
        RECT 110.740 54.125 111.120 54.505 ;
        RECT 109.320 53.465 109.700 53.845 ;
        RECT 110.740 53.465 111.120 53.845 ;
        RECT 109.320 52.805 109.700 53.185 ;
        RECT 110.740 52.805 111.120 53.185 ;
        RECT 109.320 52.145 109.700 52.525 ;
        RECT 110.740 52.145 111.120 52.525 ;
        RECT 109.320 51.485 109.700 51.865 ;
        RECT 110.740 51.485 111.120 51.865 ;
        RECT 109.320 50.825 109.700 51.205 ;
        RECT 110.740 50.825 111.120 51.205 ;
        RECT 109.320 50.165 109.700 50.545 ;
        RECT 110.740 50.165 111.120 50.545 ;
        RECT 115.225 47.805 115.605 48.185 ;
        RECT 115.885 47.805 116.265 48.185 ;
        RECT 116.545 47.805 116.925 48.185 ;
        RECT 115.225 47.145 115.605 47.525 ;
        RECT 115.885 47.145 116.265 47.525 ;
        RECT 116.545 47.145 116.925 47.525 ;
        RECT 115.225 46.485 115.605 46.865 ;
        RECT 115.885 46.485 116.265 46.865 ;
        RECT 116.545 46.485 116.925 46.865 ;
        RECT 103.530 45.105 103.910 45.485 ;
        RECT 104.190 45.105 104.570 45.485 ;
        RECT 104.850 45.105 105.230 45.485 ;
        RECT 103.530 44.445 103.910 44.825 ;
        RECT 104.190 44.445 104.570 44.825 ;
        RECT 104.850 44.445 105.230 44.825 ;
        RECT 103.530 43.785 103.910 44.165 ;
        RECT 104.190 43.785 104.570 44.165 ;
        RECT 104.850 43.785 105.230 44.165 ;
        RECT 103.530 24.905 103.910 25.285 ;
        RECT 104.190 24.905 104.570 25.285 ;
        RECT 104.850 24.905 105.230 25.285 ;
        RECT 103.530 24.245 103.910 24.625 ;
        RECT 104.190 24.245 104.570 24.625 ;
        RECT 104.850 24.245 105.230 24.625 ;
        RECT 103.530 23.585 103.910 23.965 ;
        RECT 104.190 23.585 104.570 23.965 ;
        RECT 104.850 23.585 105.230 23.965 ;
        RECT 115.225 22.205 115.605 22.585 ;
        RECT 115.885 22.205 116.265 22.585 ;
        RECT 116.545 22.205 116.925 22.585 ;
        RECT 115.225 21.545 115.605 21.925 ;
        RECT 115.885 21.545 116.265 21.925 ;
        RECT 116.545 21.545 116.925 21.925 ;
        RECT 115.225 20.885 115.605 21.265 ;
        RECT 115.885 20.885 116.265 21.265 ;
        RECT 116.545 20.885 116.925 21.265 ;
        RECT 96.980 9.100 100.945 9.150 ;
        RECT 118.975 9.150 119.500 59.890 ;
        RECT 121.030 58.745 121.410 59.125 ;
        RECT 121.030 58.085 121.410 58.465 ;
        RECT 121.030 57.425 121.410 57.805 ;
        RECT 121.030 56.765 121.410 57.145 ;
        RECT 121.030 56.105 121.410 56.485 ;
        RECT 121.030 55.445 121.410 55.825 ;
        RECT 121.030 54.785 121.410 55.165 ;
        RECT 121.030 54.125 121.410 54.505 ;
        RECT 121.030 53.465 121.410 53.845 ;
        RECT 121.030 52.805 121.410 53.185 ;
        RECT 121.030 52.145 121.410 52.525 ;
        RECT 121.030 51.485 121.410 51.865 ;
        RECT 121.030 50.825 121.410 51.205 ;
        RECT 121.030 50.165 121.410 50.545 ;
        RECT 122.415 9.150 122.940 59.890 ;
        RECT 131.315 58.745 131.695 59.125 ;
        RECT 132.735 58.745 133.115 59.125 ;
        RECT 131.315 58.085 131.695 58.465 ;
        RECT 132.735 58.085 133.115 58.465 ;
        RECT 131.315 57.425 131.695 57.805 ;
        RECT 132.735 57.425 133.115 57.805 ;
        RECT 131.315 56.765 131.695 57.145 ;
        RECT 132.735 56.765 133.115 57.145 ;
        RECT 131.315 56.105 131.695 56.485 ;
        RECT 132.735 56.105 133.115 56.485 ;
        RECT 131.315 55.445 131.695 55.825 ;
        RECT 132.735 55.445 133.115 55.825 ;
        RECT 131.315 54.785 131.695 55.165 ;
        RECT 132.735 54.785 133.115 55.165 ;
        RECT 131.315 54.125 131.695 54.505 ;
        RECT 132.735 54.125 133.115 54.505 ;
        RECT 131.315 53.465 131.695 53.845 ;
        RECT 132.735 53.465 133.115 53.845 ;
        RECT 131.315 52.805 131.695 53.185 ;
        RECT 132.735 52.805 133.115 53.185 ;
        RECT 131.315 52.145 131.695 52.525 ;
        RECT 132.735 52.145 133.115 52.525 ;
        RECT 131.315 51.485 131.695 51.865 ;
        RECT 132.735 51.485 133.115 51.865 ;
        RECT 131.315 50.825 131.695 51.205 ;
        RECT 132.735 50.825 133.115 51.205 ;
        RECT 131.315 50.165 131.695 50.545 ;
        RECT 132.735 50.165 133.115 50.545 ;
        RECT 137.220 47.805 137.600 48.185 ;
        RECT 137.880 47.805 138.260 48.185 ;
        RECT 138.540 47.805 138.920 48.185 ;
        RECT 137.220 47.145 137.600 47.525 ;
        RECT 137.880 47.145 138.260 47.525 ;
        RECT 138.540 47.145 138.920 47.525 ;
        RECT 137.220 46.485 137.600 46.865 ;
        RECT 137.880 46.485 138.260 46.865 ;
        RECT 138.540 46.485 138.920 46.865 ;
        RECT 125.525 45.105 125.905 45.485 ;
        RECT 126.185 45.105 126.565 45.485 ;
        RECT 126.845 45.105 127.225 45.485 ;
        RECT 125.525 44.445 125.905 44.825 ;
        RECT 126.185 44.445 126.565 44.825 ;
        RECT 126.845 44.445 127.225 44.825 ;
        RECT 125.525 43.785 125.905 44.165 ;
        RECT 126.185 43.785 126.565 44.165 ;
        RECT 126.845 43.785 127.225 44.165 ;
        RECT 125.525 24.905 125.905 25.285 ;
        RECT 126.185 24.905 126.565 25.285 ;
        RECT 126.845 24.905 127.225 25.285 ;
        RECT 125.525 24.245 125.905 24.625 ;
        RECT 126.185 24.245 126.565 24.625 ;
        RECT 126.845 24.245 127.225 24.625 ;
        RECT 125.525 23.585 125.905 23.965 ;
        RECT 126.185 23.585 126.565 23.965 ;
        RECT 126.845 23.585 127.225 23.965 ;
        RECT 137.220 22.205 137.600 22.585 ;
        RECT 137.880 22.205 138.260 22.585 ;
        RECT 138.540 22.205 138.920 22.585 ;
        RECT 137.220 21.545 137.600 21.925 ;
        RECT 137.880 21.545 138.260 21.925 ;
        RECT 138.540 21.545 138.920 21.925 ;
        RECT 137.220 20.885 137.600 21.265 ;
        RECT 137.880 20.885 138.260 21.265 ;
        RECT 138.540 20.885 138.920 21.265 ;
        RECT 118.975 9.100 122.940 9.150 ;
        RECT 140.970 9.150 141.495 59.890 ;
        RECT 143.025 58.745 143.405 59.125 ;
        RECT 143.025 58.085 143.405 58.465 ;
        RECT 143.025 57.425 143.405 57.805 ;
        RECT 143.025 56.765 143.405 57.145 ;
        RECT 143.025 56.105 143.405 56.485 ;
        RECT 143.025 55.445 143.405 55.825 ;
        RECT 143.025 54.785 143.405 55.165 ;
        RECT 143.025 54.125 143.405 54.505 ;
        RECT 143.025 53.465 143.405 53.845 ;
        RECT 143.025 52.805 143.405 53.185 ;
        RECT 143.025 52.145 143.405 52.525 ;
        RECT 143.025 51.485 143.405 51.865 ;
        RECT 143.025 50.825 143.405 51.205 ;
        RECT 143.025 50.165 143.405 50.545 ;
        RECT 144.410 9.150 144.935 59.890 ;
        RECT 153.310 58.745 153.690 59.125 ;
        RECT 154.730 58.745 155.110 59.125 ;
        RECT 153.310 58.085 153.690 58.465 ;
        RECT 154.730 58.085 155.110 58.465 ;
        RECT 153.310 57.425 153.690 57.805 ;
        RECT 154.730 57.425 155.110 57.805 ;
        RECT 153.310 56.765 153.690 57.145 ;
        RECT 154.730 56.765 155.110 57.145 ;
        RECT 153.310 56.105 153.690 56.485 ;
        RECT 154.730 56.105 155.110 56.485 ;
        RECT 153.310 55.445 153.690 55.825 ;
        RECT 154.730 55.445 155.110 55.825 ;
        RECT 153.310 54.785 153.690 55.165 ;
        RECT 154.730 54.785 155.110 55.165 ;
        RECT 153.310 54.125 153.690 54.505 ;
        RECT 154.730 54.125 155.110 54.505 ;
        RECT 153.310 53.465 153.690 53.845 ;
        RECT 154.730 53.465 155.110 53.845 ;
        RECT 153.310 52.805 153.690 53.185 ;
        RECT 154.730 52.805 155.110 53.185 ;
        RECT 153.310 52.145 153.690 52.525 ;
        RECT 154.730 52.145 155.110 52.525 ;
        RECT 153.310 51.485 153.690 51.865 ;
        RECT 154.730 51.485 155.110 51.865 ;
        RECT 153.310 50.825 153.690 51.205 ;
        RECT 154.730 50.825 155.110 51.205 ;
        RECT 153.310 50.165 153.690 50.545 ;
        RECT 154.730 50.165 155.110 50.545 ;
        RECT 159.215 47.805 159.595 48.185 ;
        RECT 159.875 47.805 160.255 48.185 ;
        RECT 160.535 47.805 160.915 48.185 ;
        RECT 159.215 47.145 159.595 47.525 ;
        RECT 159.875 47.145 160.255 47.525 ;
        RECT 160.535 47.145 160.915 47.525 ;
        RECT 159.215 46.485 159.595 46.865 ;
        RECT 159.875 46.485 160.255 46.865 ;
        RECT 160.535 46.485 160.915 46.865 ;
        RECT 147.520 45.105 147.900 45.485 ;
        RECT 148.180 45.105 148.560 45.485 ;
        RECT 148.840 45.105 149.220 45.485 ;
        RECT 147.520 44.445 147.900 44.825 ;
        RECT 148.180 44.445 148.560 44.825 ;
        RECT 148.840 44.445 149.220 44.825 ;
        RECT 147.520 43.785 147.900 44.165 ;
        RECT 148.180 43.785 148.560 44.165 ;
        RECT 148.840 43.785 149.220 44.165 ;
        RECT 147.520 24.905 147.900 25.285 ;
        RECT 148.180 24.905 148.560 25.285 ;
        RECT 148.840 24.905 149.220 25.285 ;
        RECT 147.520 24.245 147.900 24.625 ;
        RECT 148.180 24.245 148.560 24.625 ;
        RECT 148.840 24.245 149.220 24.625 ;
        RECT 147.520 23.585 147.900 23.965 ;
        RECT 148.180 23.585 148.560 23.965 ;
        RECT 148.840 23.585 149.220 23.965 ;
        RECT 159.215 22.205 159.595 22.585 ;
        RECT 159.875 22.205 160.255 22.585 ;
        RECT 160.535 22.205 160.915 22.585 ;
        RECT 159.215 21.545 159.595 21.925 ;
        RECT 159.875 21.545 160.255 21.925 ;
        RECT 160.535 21.545 160.915 21.925 ;
        RECT 159.215 20.885 159.595 21.265 ;
        RECT 159.875 20.885 160.255 21.265 ;
        RECT 160.535 20.885 160.915 21.265 ;
        RECT 140.970 9.100 144.935 9.150 ;
        RECT 162.965 9.150 163.490 59.890 ;
        RECT 165.020 58.745 165.400 59.125 ;
        RECT 165.020 58.085 165.400 58.465 ;
        RECT 165.020 57.425 165.400 57.805 ;
        RECT 165.020 56.765 165.400 57.145 ;
        RECT 165.020 56.105 165.400 56.485 ;
        RECT 165.020 55.445 165.400 55.825 ;
        RECT 165.020 54.785 165.400 55.165 ;
        RECT 165.020 54.125 165.400 54.505 ;
        RECT 165.020 53.465 165.400 53.845 ;
        RECT 165.020 52.805 165.400 53.185 ;
        RECT 165.020 52.145 165.400 52.525 ;
        RECT 165.020 51.485 165.400 51.865 ;
        RECT 165.020 50.825 165.400 51.205 ;
        RECT 165.020 50.165 165.400 50.545 ;
        RECT 166.405 9.150 166.930 59.890 ;
        RECT 175.305 58.745 175.685 59.125 ;
        RECT 175.305 58.085 175.685 58.465 ;
        RECT 175.305 57.425 175.685 57.805 ;
        RECT 175.305 56.765 175.685 57.145 ;
        RECT 175.305 56.105 175.685 56.485 ;
        RECT 175.305 55.445 175.685 55.825 ;
        RECT 175.305 54.785 175.685 55.165 ;
        RECT 177.150 55.115 177.530 55.495 ;
        RECT 178.935 55.115 179.315 55.495 ;
        RECT 181.790 55.115 182.170 55.495 ;
        RECT 183.575 55.115 183.955 55.495 ;
        RECT 186.430 55.115 186.810 55.495 ;
        RECT 188.215 55.115 188.595 55.495 ;
        RECT 191.070 55.115 191.450 55.495 ;
        RECT 192.855 55.115 193.235 55.495 ;
        RECT 175.305 54.125 175.685 54.505 ;
        RECT 177.150 54.455 177.530 54.835 ;
        RECT 178.935 54.455 179.315 54.835 ;
        RECT 181.790 54.455 182.170 54.835 ;
        RECT 183.575 54.455 183.955 54.835 ;
        RECT 186.430 54.455 186.810 54.835 ;
        RECT 188.215 54.455 188.595 54.835 ;
        RECT 191.070 54.455 191.450 54.835 ;
        RECT 192.855 54.455 193.235 54.835 ;
        RECT 175.305 53.465 175.685 53.845 ;
        RECT 177.150 53.795 177.530 54.175 ;
        RECT 178.935 53.795 179.315 54.175 ;
        RECT 181.790 53.795 182.170 54.175 ;
        RECT 183.575 53.795 183.955 54.175 ;
        RECT 186.430 53.795 186.810 54.175 ;
        RECT 188.215 53.795 188.595 54.175 ;
        RECT 191.070 53.795 191.450 54.175 ;
        RECT 192.855 53.795 193.235 54.175 ;
        RECT 175.305 52.805 175.685 53.185 ;
        RECT 177.150 53.135 177.530 53.515 ;
        RECT 178.935 53.135 179.315 53.515 ;
        RECT 181.790 53.135 182.170 53.515 ;
        RECT 183.575 53.135 183.955 53.515 ;
        RECT 186.430 53.135 186.810 53.515 ;
        RECT 188.215 53.135 188.595 53.515 ;
        RECT 191.070 53.135 191.450 53.515 ;
        RECT 192.855 53.135 193.235 53.515 ;
        RECT 175.305 52.145 175.685 52.525 ;
        RECT 177.150 52.475 177.530 52.855 ;
        RECT 178.935 52.475 179.315 52.855 ;
        RECT 181.790 52.475 182.170 52.855 ;
        RECT 183.575 52.475 183.955 52.855 ;
        RECT 186.430 52.475 186.810 52.855 ;
        RECT 188.215 52.475 188.595 52.855 ;
        RECT 191.070 52.475 191.450 52.855 ;
        RECT 192.855 52.475 193.235 52.855 ;
        RECT 175.305 51.485 175.685 51.865 ;
        RECT 177.150 51.815 177.530 52.195 ;
        RECT 178.935 51.815 179.315 52.195 ;
        RECT 181.790 51.815 182.170 52.195 ;
        RECT 183.575 51.815 183.955 52.195 ;
        RECT 186.430 51.815 186.810 52.195 ;
        RECT 188.215 51.815 188.595 52.195 ;
        RECT 191.070 51.815 191.450 52.195 ;
        RECT 192.855 51.815 193.235 52.195 ;
        RECT 175.305 50.825 175.685 51.205 ;
        RECT 177.150 51.155 177.530 51.535 ;
        RECT 178.935 51.155 179.315 51.535 ;
        RECT 181.790 51.155 182.170 51.535 ;
        RECT 183.575 51.155 183.955 51.535 ;
        RECT 186.430 51.155 186.810 51.535 ;
        RECT 188.215 51.155 188.595 51.535 ;
        RECT 191.070 51.155 191.450 51.535 ;
        RECT 192.855 51.155 193.235 51.535 ;
        RECT 175.305 50.165 175.685 50.545 ;
        RECT 177.150 50.495 177.530 50.875 ;
        RECT 178.935 50.495 179.315 50.875 ;
        RECT 181.790 50.495 182.170 50.875 ;
        RECT 183.575 50.495 183.955 50.875 ;
        RECT 186.430 50.495 186.810 50.875 ;
        RECT 188.215 50.495 188.595 50.875 ;
        RECT 191.070 50.495 191.450 50.875 ;
        RECT 192.855 50.495 193.235 50.875 ;
        RECT 177.910 47.805 178.290 48.185 ;
        RECT 177.910 47.145 178.290 47.525 ;
        RECT 177.910 46.485 178.290 46.865 ;
        RECT 169.515 45.105 169.895 45.485 ;
        RECT 170.175 45.105 170.555 45.485 ;
        RECT 170.835 45.105 171.215 45.485 ;
        RECT 191.830 45.105 192.210 45.485 ;
        RECT 169.515 44.445 169.895 44.825 ;
        RECT 170.175 44.445 170.555 44.825 ;
        RECT 170.835 44.445 171.215 44.825 ;
        RECT 191.830 44.445 192.210 44.825 ;
        RECT 169.515 43.785 169.895 44.165 ;
        RECT 170.175 43.785 170.555 44.165 ;
        RECT 170.835 43.785 171.215 44.165 ;
        RECT 191.830 43.785 192.210 44.165 ;
        RECT 169.515 24.905 169.895 25.285 ;
        RECT 170.175 24.905 170.555 25.285 ;
        RECT 170.835 24.905 171.215 25.285 ;
        RECT 187.190 24.905 187.570 25.285 ;
        RECT 169.515 24.245 169.895 24.625 ;
        RECT 170.175 24.245 170.555 24.625 ;
        RECT 170.835 24.245 171.215 24.625 ;
        RECT 187.190 24.245 187.570 24.625 ;
        RECT 169.515 23.585 169.895 23.965 ;
        RECT 170.175 23.585 170.555 23.965 ;
        RECT 170.835 23.585 171.215 23.965 ;
        RECT 187.190 23.585 187.570 23.965 ;
        RECT 182.550 22.205 182.930 22.585 ;
        RECT 182.550 21.545 182.930 21.925 ;
        RECT 182.550 20.885 182.930 21.265 ;
        RECT 177.150 18.115 177.530 18.495 ;
        RECT 178.935 18.115 179.315 18.495 ;
        RECT 181.790 18.115 182.170 18.495 ;
        RECT 183.575 18.115 183.955 18.495 ;
        RECT 186.430 18.115 186.810 18.495 ;
        RECT 188.215 18.115 188.595 18.495 ;
        RECT 191.070 18.115 191.450 18.495 ;
        RECT 192.855 18.115 193.235 18.495 ;
        RECT 177.150 17.455 177.530 17.835 ;
        RECT 178.935 17.455 179.315 17.835 ;
        RECT 181.790 17.455 182.170 17.835 ;
        RECT 183.575 17.455 183.955 17.835 ;
        RECT 186.430 17.455 186.810 17.835 ;
        RECT 188.215 17.455 188.595 17.835 ;
        RECT 191.070 17.455 191.450 17.835 ;
        RECT 192.855 17.455 193.235 17.835 ;
        RECT 177.150 16.795 177.530 17.175 ;
        RECT 178.935 16.795 179.315 17.175 ;
        RECT 181.790 16.795 182.170 17.175 ;
        RECT 183.575 16.795 183.955 17.175 ;
        RECT 186.430 16.795 186.810 17.175 ;
        RECT 188.215 16.795 188.595 17.175 ;
        RECT 191.070 16.795 191.450 17.175 ;
        RECT 192.855 16.795 193.235 17.175 ;
        RECT 177.150 16.135 177.530 16.515 ;
        RECT 178.935 16.135 179.315 16.515 ;
        RECT 181.790 16.135 182.170 16.515 ;
        RECT 183.575 16.135 183.955 16.515 ;
        RECT 186.430 16.135 186.810 16.515 ;
        RECT 188.215 16.135 188.595 16.515 ;
        RECT 191.070 16.135 191.450 16.515 ;
        RECT 192.855 16.135 193.235 16.515 ;
        RECT 177.150 15.475 177.530 15.855 ;
        RECT 178.935 15.475 179.315 15.855 ;
        RECT 181.790 15.475 182.170 15.855 ;
        RECT 183.575 15.475 183.955 15.855 ;
        RECT 186.430 15.475 186.810 15.855 ;
        RECT 188.215 15.475 188.595 15.855 ;
        RECT 191.070 15.475 191.450 15.855 ;
        RECT 192.855 15.475 193.235 15.855 ;
        RECT 177.150 14.815 177.530 15.195 ;
        RECT 178.935 14.815 179.315 15.195 ;
        RECT 181.790 14.815 182.170 15.195 ;
        RECT 183.575 14.815 183.955 15.195 ;
        RECT 186.430 14.815 186.810 15.195 ;
        RECT 188.215 14.815 188.595 15.195 ;
        RECT 191.070 14.815 191.450 15.195 ;
        RECT 192.855 14.815 193.235 15.195 ;
        RECT 177.150 14.155 177.530 14.535 ;
        RECT 178.935 14.155 179.315 14.535 ;
        RECT 181.790 14.155 182.170 14.535 ;
        RECT 183.575 14.155 183.955 14.535 ;
        RECT 186.430 14.155 186.810 14.535 ;
        RECT 188.215 14.155 188.595 14.535 ;
        RECT 191.070 14.155 191.450 14.535 ;
        RECT 192.855 14.155 193.235 14.535 ;
        RECT 177.150 13.495 177.530 13.875 ;
        RECT 178.935 13.495 179.315 13.875 ;
        RECT 181.790 13.495 182.170 13.875 ;
        RECT 183.575 13.495 183.955 13.875 ;
        RECT 186.430 13.495 186.810 13.875 ;
        RECT 188.215 13.495 188.595 13.875 ;
        RECT 191.070 13.495 191.450 13.875 ;
        RECT 192.855 13.495 193.235 13.875 ;
        RECT 177.150 12.835 177.530 13.215 ;
        RECT 178.935 12.835 179.315 13.215 ;
        RECT 181.790 12.835 182.170 13.215 ;
        RECT 183.575 12.835 183.955 13.215 ;
        RECT 186.430 12.835 186.810 13.215 ;
        RECT 188.215 12.835 188.595 13.215 ;
        RECT 191.070 12.835 191.450 13.215 ;
        RECT 192.855 12.835 193.235 13.215 ;
        RECT 177.150 12.175 177.530 12.555 ;
        RECT 178.935 12.175 179.315 12.555 ;
        RECT 181.790 12.175 182.170 12.555 ;
        RECT 183.575 12.175 183.955 12.555 ;
        RECT 186.430 12.175 186.810 12.555 ;
        RECT 188.215 12.175 188.595 12.555 ;
        RECT 191.070 12.175 191.450 12.555 ;
        RECT 192.855 12.175 193.235 12.555 ;
        RECT 177.150 11.515 177.530 11.895 ;
        RECT 178.935 11.515 179.315 11.895 ;
        RECT 181.790 11.515 182.170 11.895 ;
        RECT 183.575 11.515 183.955 11.895 ;
        RECT 186.430 11.515 186.810 11.895 ;
        RECT 188.215 11.515 188.595 11.895 ;
        RECT 191.070 11.515 191.450 11.895 ;
        RECT 192.855 11.515 193.235 11.895 ;
        RECT 177.150 10.855 177.530 11.235 ;
        RECT 178.935 10.855 179.315 11.235 ;
        RECT 181.790 10.855 182.170 11.235 ;
        RECT 183.575 10.855 183.955 11.235 ;
        RECT 186.430 10.855 186.810 11.235 ;
        RECT 188.215 10.855 188.595 11.235 ;
        RECT 191.070 10.855 191.450 11.235 ;
        RECT 192.855 10.855 193.235 11.235 ;
        RECT 177.150 10.195 177.530 10.575 ;
        RECT 178.935 10.195 179.315 10.575 ;
        RECT 181.790 10.195 182.170 10.575 ;
        RECT 183.575 10.195 183.955 10.575 ;
        RECT 186.430 10.195 186.810 10.575 ;
        RECT 188.215 10.195 188.595 10.575 ;
        RECT 191.070 10.195 191.450 10.575 ;
        RECT 192.855 10.195 193.235 10.575 ;
        RECT 177.150 9.535 177.530 9.915 ;
        RECT 178.935 9.535 179.315 9.915 ;
        RECT 181.790 9.535 182.170 9.915 ;
        RECT 183.575 9.535 183.955 9.915 ;
        RECT 186.430 9.535 186.810 9.915 ;
        RECT 188.215 9.535 188.595 9.915 ;
        RECT 191.070 9.535 191.450 9.915 ;
        RECT 192.855 9.535 193.235 9.915 ;
        RECT 162.965 9.100 166.930 9.150 ;
        RECT 9.000 8.770 20.385 9.100 ;
        RECT 9.000 8.750 12.965 8.770 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 0.850 4.690 1.230 5.070 ;
        RECT 1.990 4.690 2.370 5.070 ;
        RECT 8.030 4.720 8.410 5.100 ;
        RECT 8.690 4.720 9.070 5.100 ;
        RECT 9.350 4.720 9.730 5.100 ;
        RECT 14.560 4.690 14.940 5.070 ;
        RECT 15.220 4.690 15.600 5.070 ;
        RECT 15.880 4.690 16.260 5.070 ;
        RECT 17.920 4.690 18.300 5.070 ;
        RECT 18.580 4.690 18.960 5.070 ;
        RECT 19.240 4.690 19.620 5.070 ;
        RECT 3.490 2.950 3.860 4.550 ;
        RECT 20.055 4.150 20.385 8.770 ;
        RECT 30.995 8.770 38.575 9.100 ;
        RECT 30.995 8.750 34.960 8.770 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 26.220 4.720 26.600 5.100 ;
        RECT 26.880 4.720 27.260 5.100 ;
        RECT 27.540 4.720 27.920 5.100 ;
        RECT 32.750 4.690 33.130 5.070 ;
        RECT 33.410 4.690 33.790 5.070 ;
        RECT 34.070 4.690 34.450 5.070 ;
        RECT 36.110 4.690 36.490 5.070 ;
        RECT 36.770 4.690 37.150 5.070 ;
        RECT 37.430 4.690 37.810 5.070 ;
        RECT 4.170 3.420 4.550 3.800 ;
        RECT 20.030 3.770 20.410 4.150 ;
        RECT 3.490 2.580 4.190 2.950 ;
        RECT 4.580 2.760 4.960 3.140 ;
        RECT 6.995 2.950 10.205 3.300 ;
        RECT 3.820 2.305 4.190 2.580 ;
        RECT 6.995 2.305 7.345 2.950 ;
        RECT 11.480 2.760 13.000 3.255 ;
        RECT 14.945 3.125 15.325 3.150 ;
        RECT 13.865 2.795 15.325 3.125 ;
        RECT 11.480 2.600 11.890 2.760 ;
        RECT 3.820 1.955 7.345 2.305 ;
        RECT 7.645 2.250 11.890 2.600 ;
        RECT 12.090 1.885 12.470 1.910 ;
        RECT 13.865 1.885 14.195 2.795 ;
        RECT 14.945 2.770 15.325 2.795 ;
        RECT 21.680 2.950 22.050 4.550 ;
        RECT 38.245 4.150 38.575 8.770 ;
        RECT 52.990 8.770 72.715 9.100 ;
        RECT 52.990 8.750 56.955 8.770 ;
        RECT 42.110 8.090 42.490 8.470 ;
        RECT 56.940 8.090 57.320 8.470 ;
        RECT 42.110 7.430 42.490 7.810 ;
        RECT 56.940 7.430 57.320 7.810 ;
        RECT 42.110 6.770 42.490 7.150 ;
        RECT 56.940 6.770 57.320 7.150 ;
        RECT 39.490 4.690 39.870 5.070 ;
        RECT 45.530 4.720 45.910 5.100 ;
        RECT 46.190 4.720 46.570 5.100 ;
        RECT 46.850 4.720 47.230 5.100 ;
        RECT 52.060 4.690 52.440 5.070 ;
        RECT 52.720 4.690 53.100 5.070 ;
        RECT 53.380 4.690 53.760 5.070 ;
        RECT 60.360 4.720 60.740 5.100 ;
        RECT 61.020 4.720 61.400 5.100 ;
        RECT 61.680 4.720 62.060 5.100 ;
        RECT 66.890 4.690 67.270 5.070 ;
        RECT 67.550 4.690 67.930 5.070 ;
        RECT 68.210 4.690 68.590 5.070 ;
        RECT 70.250 4.690 70.630 5.070 ;
        RECT 70.910 4.690 71.290 5.070 ;
        RECT 71.570 4.690 71.950 5.070 ;
        RECT 22.360 3.420 22.740 3.800 ;
        RECT 38.220 3.770 38.600 4.150 ;
        RECT 21.680 2.580 22.380 2.950 ;
        RECT 22.770 2.760 23.150 3.140 ;
        RECT 25.185 2.950 28.395 3.300 ;
        RECT 22.010 2.305 22.380 2.580 ;
        RECT 25.185 2.305 25.535 2.950 ;
        RECT 29.670 2.760 31.190 3.255 ;
        RECT 33.135 3.125 33.515 3.150 ;
        RECT 32.055 2.795 33.515 3.125 ;
        RECT 29.670 2.600 30.080 2.760 ;
        RECT 22.010 1.955 25.535 2.305 ;
        RECT 25.835 2.250 30.080 2.600 ;
        RECT 12.090 1.555 14.195 1.885 ;
        RECT 30.280 1.885 30.660 1.910 ;
        RECT 32.055 1.885 32.385 2.795 ;
        RECT 33.135 2.770 33.515 2.795 ;
        RECT 40.990 2.950 41.360 4.550 ;
        RECT 41.670 3.420 42.050 3.800 ;
        RECT 40.990 2.580 41.690 2.950 ;
        RECT 42.080 2.760 42.460 3.140 ;
        RECT 44.495 2.950 47.705 3.300 ;
        RECT 41.320 2.305 41.690 2.580 ;
        RECT 44.495 2.305 44.845 2.950 ;
        RECT 48.980 2.760 50.500 3.255 ;
        RECT 52.445 3.125 52.825 3.150 ;
        RECT 51.365 2.795 52.825 3.125 ;
        RECT 48.980 2.600 49.390 2.760 ;
        RECT 41.320 1.955 44.845 2.305 ;
        RECT 45.145 2.250 49.390 2.600 ;
        RECT 30.280 1.555 32.385 1.885 ;
        RECT 49.590 1.885 49.970 1.910 ;
        RECT 51.365 1.885 51.695 2.795 ;
        RECT 52.445 2.770 52.825 2.795 ;
        RECT 55.820 2.950 56.190 4.550 ;
        RECT 72.385 4.150 72.715 8.770 ;
        RECT 74.985 8.770 81.675 9.100 ;
        RECT 74.985 8.750 78.950 8.770 ;
        RECT 73.630 4.690 74.010 5.070 ;
        RECT 74.630 4.690 75.010 5.070 ;
        RECT 75.290 4.690 75.670 5.070 ;
        RECT 75.950 4.690 76.330 5.070 ;
        RECT 76.870 4.690 77.250 5.070 ;
        RECT 77.530 4.690 77.910 5.070 ;
        RECT 78.190 4.690 78.570 5.070 ;
        RECT 79.210 4.690 79.590 5.070 ;
        RECT 79.870 4.690 80.250 5.070 ;
        RECT 80.530 4.690 80.910 5.070 ;
        RECT 81.345 4.150 81.675 8.770 ;
        RECT 96.980 8.770 104.075 9.100 ;
        RECT 96.980 8.750 100.945 8.770 ;
        RECT 82.470 4.690 82.850 5.070 ;
        RECT 83.130 4.690 83.510 5.070 ;
        RECT 83.790 4.690 84.170 5.070 ;
        RECT 84.710 4.690 85.090 5.070 ;
        RECT 85.370 4.690 85.750 5.070 ;
        RECT 86.030 4.690 86.410 5.070 ;
        RECT 86.950 4.690 87.330 5.070 ;
        RECT 87.610 4.690 87.990 5.070 ;
        RECT 88.270 4.690 88.650 5.070 ;
        RECT 89.190 4.690 89.570 5.070 ;
        RECT 89.850 4.690 90.230 5.070 ;
        RECT 90.510 4.690 90.890 5.070 ;
        RECT 91.430 4.690 91.810 5.070 ;
        RECT 92.090 4.690 92.470 5.070 ;
        RECT 92.750 4.690 93.130 5.070 ;
        RECT 93.790 4.690 94.170 5.070 ;
        RECT 94.790 4.690 95.170 5.070 ;
        RECT 95.450 4.690 95.830 5.070 ;
        RECT 96.110 4.690 96.490 5.070 ;
        RECT 97.030 4.690 97.410 5.070 ;
        RECT 97.690 4.690 98.070 5.070 ;
        RECT 98.350 4.690 98.730 5.070 ;
        RECT 99.270 4.690 99.650 5.070 ;
        RECT 99.930 4.690 100.310 5.070 ;
        RECT 100.590 4.690 100.970 5.070 ;
        RECT 101.610 4.690 101.990 5.070 ;
        RECT 102.270 4.690 102.650 5.070 ;
        RECT 102.930 4.690 103.310 5.070 ;
        RECT 103.745 4.150 104.075 8.770 ;
        RECT 118.975 8.770 124.235 9.100 ;
        RECT 118.975 8.750 122.940 8.770 ;
        RECT 104.870 4.690 105.250 5.070 ;
        RECT 105.530 4.690 105.910 5.070 ;
        RECT 106.190 4.690 106.570 5.070 ;
        RECT 107.110 4.690 107.490 5.070 ;
        RECT 107.770 4.690 108.150 5.070 ;
        RECT 108.430 4.690 108.810 5.070 ;
        RECT 109.350 4.690 109.730 5.070 ;
        RECT 110.010 4.690 110.390 5.070 ;
        RECT 110.670 4.690 111.050 5.070 ;
        RECT 111.590 4.690 111.970 5.070 ;
        RECT 112.250 4.690 112.630 5.070 ;
        RECT 112.910 4.690 113.290 5.070 ;
        RECT 113.950 4.690 114.330 5.070 ;
        RECT 114.950 4.690 115.330 5.070 ;
        RECT 115.610 4.690 115.990 5.070 ;
        RECT 116.270 4.690 116.650 5.070 ;
        RECT 117.190 4.690 117.570 5.070 ;
        RECT 117.850 4.690 118.230 5.070 ;
        RECT 118.510 4.690 118.890 5.070 ;
        RECT 119.430 4.690 119.810 5.070 ;
        RECT 120.090 4.690 120.470 5.070 ;
        RECT 120.750 4.690 121.130 5.070 ;
        RECT 121.770 4.690 122.150 5.070 ;
        RECT 122.430 4.690 122.810 5.070 ;
        RECT 123.090 4.690 123.470 5.070 ;
        RECT 123.905 4.150 124.235 8.770 ;
        RECT 140.970 8.770 146.635 9.100 ;
        RECT 140.970 8.750 144.935 8.770 ;
        RECT 125.030 4.690 125.410 5.070 ;
        RECT 125.690 4.690 126.070 5.070 ;
        RECT 126.350 4.690 126.730 5.070 ;
        RECT 127.270 4.690 127.650 5.070 ;
        RECT 127.930 4.690 128.310 5.070 ;
        RECT 128.590 4.690 128.970 5.070 ;
        RECT 129.510 4.690 129.890 5.070 ;
        RECT 130.170 4.690 130.550 5.070 ;
        RECT 130.830 4.690 131.210 5.070 ;
        RECT 131.750 4.690 132.130 5.070 ;
        RECT 132.410 4.690 132.790 5.070 ;
        RECT 133.070 4.690 133.450 5.070 ;
        RECT 134.110 4.690 134.490 5.070 ;
        RECT 135.110 4.690 135.490 5.070 ;
        RECT 135.770 4.690 136.150 5.070 ;
        RECT 136.430 4.690 136.810 5.070 ;
        RECT 137.350 4.690 137.730 5.070 ;
        RECT 138.010 4.690 138.390 5.070 ;
        RECT 138.670 4.690 139.050 5.070 ;
        RECT 139.590 4.690 139.970 5.070 ;
        RECT 140.250 4.690 140.630 5.070 ;
        RECT 140.910 4.690 141.290 5.070 ;
        RECT 141.830 4.690 142.210 5.070 ;
        RECT 142.490 4.690 142.870 5.070 ;
        RECT 143.150 4.690 143.530 5.070 ;
        RECT 144.170 4.690 144.550 5.070 ;
        RECT 144.830 4.690 145.210 5.070 ;
        RECT 145.490 4.690 145.870 5.070 ;
        RECT 146.305 4.150 146.635 8.770 ;
        RECT 162.965 8.770 169.035 9.100 ;
        RECT 177.150 8.875 177.530 9.255 ;
        RECT 178.935 8.875 179.315 9.255 ;
        RECT 181.790 8.875 182.170 9.255 ;
        RECT 183.575 8.875 183.955 9.255 ;
        RECT 186.430 8.875 186.810 9.255 ;
        RECT 188.215 8.875 188.595 9.255 ;
        RECT 191.070 8.875 191.450 9.255 ;
        RECT 192.855 8.875 193.235 9.255 ;
        RECT 162.965 8.750 166.930 8.770 ;
        RECT 147.430 4.690 147.810 5.070 ;
        RECT 148.090 4.690 148.470 5.070 ;
        RECT 148.750 4.690 149.130 5.070 ;
        RECT 149.670 4.690 150.050 5.070 ;
        RECT 150.330 4.690 150.710 5.070 ;
        RECT 150.990 4.690 151.370 5.070 ;
        RECT 151.910 4.690 152.290 5.070 ;
        RECT 152.570 4.690 152.950 5.070 ;
        RECT 153.230 4.690 153.610 5.070 ;
        RECT 154.270 4.690 154.650 5.070 ;
        RECT 155.270 4.690 155.650 5.070 ;
        RECT 155.930 4.690 156.310 5.070 ;
        RECT 156.590 4.690 156.970 5.070 ;
        RECT 157.510 4.690 157.890 5.070 ;
        RECT 158.170 4.690 158.550 5.070 ;
        RECT 158.830 4.690 159.210 5.070 ;
        RECT 159.750 4.690 160.130 5.070 ;
        RECT 160.410 4.690 160.790 5.070 ;
        RECT 161.070 4.690 161.450 5.070 ;
        RECT 161.990 4.690 162.370 5.070 ;
        RECT 162.650 4.690 163.030 5.070 ;
        RECT 163.310 4.690 163.690 5.070 ;
        RECT 164.230 4.690 164.610 5.070 ;
        RECT 164.890 4.690 165.270 5.070 ;
        RECT 165.550 4.690 165.930 5.070 ;
        RECT 166.570 4.690 166.950 5.070 ;
        RECT 167.230 4.690 167.610 5.070 ;
        RECT 167.890 4.690 168.270 5.070 ;
        RECT 168.705 4.150 169.035 8.770 ;
        RECT 169.830 4.690 170.210 5.070 ;
        RECT 170.490 4.690 170.870 5.070 ;
        RECT 171.150 4.690 171.530 5.070 ;
        RECT 172.070 4.690 172.450 5.070 ;
        RECT 172.730 4.690 173.110 5.070 ;
        RECT 173.390 4.690 173.770 5.070 ;
        RECT 174.410 4.690 174.790 5.070 ;
        RECT 56.500 3.420 56.880 3.800 ;
        RECT 72.360 3.770 72.740 4.150 ;
        RECT 81.320 3.770 81.700 4.150 ;
        RECT 103.720 3.770 104.100 4.150 ;
        RECT 123.880 3.770 124.260 4.150 ;
        RECT 146.280 3.770 146.660 4.150 ;
        RECT 168.680 3.770 169.060 4.150 ;
        RECT 55.820 2.580 56.520 2.950 ;
        RECT 56.910 2.760 57.290 3.140 ;
        RECT 59.325 2.950 62.535 3.300 ;
        RECT 56.150 2.305 56.520 2.580 ;
        RECT 59.325 2.305 59.675 2.950 ;
        RECT 63.810 2.760 65.330 3.255 ;
        RECT 67.275 3.125 67.655 3.150 ;
        RECT 66.195 2.795 67.655 3.125 ;
        RECT 63.810 2.600 64.220 2.760 ;
        RECT 56.150 1.955 59.675 2.305 ;
        RECT 59.975 2.250 64.220 2.600 ;
        RECT 49.590 1.555 51.695 1.885 ;
        RECT 64.420 1.885 64.800 1.910 ;
        RECT 66.195 1.885 66.525 2.795 ;
        RECT 67.275 2.770 67.655 2.795 ;
        RECT 64.420 1.555 66.525 1.885 ;
        RECT 12.090 1.530 12.470 1.555 ;
        RECT 30.280 1.530 30.660 1.555 ;
        RECT 49.590 1.530 49.970 1.555 ;
        RECT 64.420 1.530 64.800 1.555 ;
        RECT 0.850 0.770 1.230 1.150 ;
        RECT 1.990 0.770 2.370 1.150 ;
        RECT 7.430 0.770 7.810 1.150 ;
        RECT 8.090 0.770 8.470 1.150 ;
        RECT 8.750 0.770 9.130 1.150 ;
        RECT 14.300 0.770 14.680 1.150 ;
        RECT 15.620 0.770 16.000 1.150 ;
        RECT 17.660 0.770 18.040 1.150 ;
        RECT 18.980 0.770 19.360 1.150 ;
        RECT 25.620 0.770 26.000 1.150 ;
        RECT 26.280 0.770 26.660 1.150 ;
        RECT 26.940 0.770 27.320 1.150 ;
        RECT 32.490 0.770 32.870 1.150 ;
        RECT 33.810 0.770 34.190 1.150 ;
        RECT 35.850 0.770 36.230 1.150 ;
        RECT 37.170 0.770 37.550 1.150 ;
        RECT 39.490 0.770 39.870 1.150 ;
        RECT 44.930 0.770 45.310 1.150 ;
        RECT 45.590 0.770 45.970 1.150 ;
        RECT 46.250 0.770 46.630 1.150 ;
        RECT 51.800 0.770 52.180 1.150 ;
        RECT 53.120 0.770 53.500 1.150 ;
        RECT 59.760 0.770 60.140 1.150 ;
        RECT 60.420 0.770 60.800 1.150 ;
        RECT 61.080 0.770 61.460 1.150 ;
        RECT 66.630 0.770 67.010 1.150 ;
        RECT 67.950 0.770 68.330 1.150 ;
        RECT 69.990 0.770 70.370 1.150 ;
        RECT 71.310 0.770 71.690 1.150 ;
        RECT 73.630 0.770 74.010 1.150 ;
        RECT 74.630 0.770 75.010 1.150 ;
        RECT 75.290 0.770 75.670 1.150 ;
        RECT 75.950 0.770 76.330 1.150 ;
        RECT 76.870 0.770 77.250 1.150 ;
        RECT 77.530 0.770 77.910 1.150 ;
        RECT 78.190 0.770 78.570 1.150 ;
        RECT 78.950 0.770 79.330 1.150 ;
        RECT 80.270 0.770 80.650 1.150 ;
        RECT 82.470 0.770 82.850 1.150 ;
        RECT 83.130 0.770 83.510 1.150 ;
        RECT 83.790 0.770 84.170 1.150 ;
        RECT 84.710 0.770 85.090 1.150 ;
        RECT 85.370 0.770 85.750 1.150 ;
        RECT 86.030 0.770 86.410 1.150 ;
        RECT 86.950 0.770 87.330 1.150 ;
        RECT 87.610 0.770 87.990 1.150 ;
        RECT 88.270 0.770 88.650 1.150 ;
        RECT 89.190 0.770 89.570 1.150 ;
        RECT 89.850 0.770 90.230 1.150 ;
        RECT 90.510 0.770 90.890 1.150 ;
        RECT 91.430 0.770 91.810 1.150 ;
        RECT 92.090 0.770 92.470 1.150 ;
        RECT 92.750 0.770 93.130 1.150 ;
        RECT 93.790 0.770 94.170 1.150 ;
        RECT 94.790 0.770 95.170 1.150 ;
        RECT 95.450 0.770 95.830 1.150 ;
        RECT 96.110 0.770 96.490 1.150 ;
        RECT 97.030 0.770 97.410 1.150 ;
        RECT 97.690 0.770 98.070 1.150 ;
        RECT 98.350 0.770 98.730 1.150 ;
        RECT 99.270 0.770 99.650 1.150 ;
        RECT 99.930 0.770 100.310 1.150 ;
        RECT 100.590 0.770 100.970 1.150 ;
        RECT 101.350 0.770 101.730 1.150 ;
        RECT 102.670 0.770 103.050 1.150 ;
        RECT 104.870 0.770 105.250 1.150 ;
        RECT 105.530 0.770 105.910 1.150 ;
        RECT 106.190 0.770 106.570 1.150 ;
        RECT 107.110 0.770 107.490 1.150 ;
        RECT 107.770 0.770 108.150 1.150 ;
        RECT 108.430 0.770 108.810 1.150 ;
        RECT 109.350 0.770 109.730 1.150 ;
        RECT 110.010 0.770 110.390 1.150 ;
        RECT 110.670 0.770 111.050 1.150 ;
        RECT 111.590 0.770 111.970 1.150 ;
        RECT 112.250 0.770 112.630 1.150 ;
        RECT 112.910 0.770 113.290 1.150 ;
        RECT 113.950 0.770 114.330 1.150 ;
        RECT 114.950 0.770 115.330 1.150 ;
        RECT 115.610 0.770 115.990 1.150 ;
        RECT 116.270 0.770 116.650 1.150 ;
        RECT 117.190 0.770 117.570 1.150 ;
        RECT 117.850 0.770 118.230 1.150 ;
        RECT 118.510 0.770 118.890 1.150 ;
        RECT 119.430 0.770 119.810 1.150 ;
        RECT 120.090 0.770 120.470 1.150 ;
        RECT 120.750 0.770 121.130 1.150 ;
        RECT 121.510 0.770 121.890 1.150 ;
        RECT 122.830 0.770 123.210 1.150 ;
        RECT 125.030 0.770 125.410 1.150 ;
        RECT 125.690 0.770 126.070 1.150 ;
        RECT 126.350 0.770 126.730 1.150 ;
        RECT 127.270 0.770 127.650 1.150 ;
        RECT 127.930 0.770 128.310 1.150 ;
        RECT 128.590 0.770 128.970 1.150 ;
        RECT 129.510 0.770 129.890 1.150 ;
        RECT 130.170 0.770 130.550 1.150 ;
        RECT 130.830 0.770 131.210 1.150 ;
        RECT 131.750 0.770 132.130 1.150 ;
        RECT 132.410 0.770 132.790 1.150 ;
        RECT 133.070 0.770 133.450 1.150 ;
        RECT 134.110 0.770 134.490 1.150 ;
        RECT 135.110 0.770 135.490 1.150 ;
        RECT 135.770 0.770 136.150 1.150 ;
        RECT 136.430 0.770 136.810 1.150 ;
        RECT 137.350 0.770 137.730 1.150 ;
        RECT 138.010 0.770 138.390 1.150 ;
        RECT 138.670 0.770 139.050 1.150 ;
        RECT 139.590 0.770 139.970 1.150 ;
        RECT 140.250 0.770 140.630 1.150 ;
        RECT 140.910 0.770 141.290 1.150 ;
        RECT 141.830 0.770 142.210 1.150 ;
        RECT 142.490 0.770 142.870 1.150 ;
        RECT 143.150 0.770 143.530 1.150 ;
        RECT 143.910 0.770 144.290 1.150 ;
        RECT 145.230 0.770 145.610 1.150 ;
        RECT 147.430 0.770 147.810 1.150 ;
        RECT 148.090 0.770 148.470 1.150 ;
        RECT 148.750 0.770 149.130 1.150 ;
        RECT 149.670 0.770 150.050 1.150 ;
        RECT 150.330 0.770 150.710 1.150 ;
        RECT 150.990 0.770 151.370 1.150 ;
        RECT 151.910 0.770 152.290 1.150 ;
        RECT 152.570 0.770 152.950 1.150 ;
        RECT 153.230 0.770 153.610 1.150 ;
        RECT 154.270 0.770 154.650 1.150 ;
        RECT 155.270 0.770 155.650 1.150 ;
        RECT 155.930 0.770 156.310 1.150 ;
        RECT 156.590 0.770 156.970 1.150 ;
        RECT 157.510 0.770 157.890 1.150 ;
        RECT 158.170 0.770 158.550 1.150 ;
        RECT 158.830 0.770 159.210 1.150 ;
        RECT 159.750 0.770 160.130 1.150 ;
        RECT 160.410 0.770 160.790 1.150 ;
        RECT 161.070 0.770 161.450 1.150 ;
        RECT 161.990 0.770 162.370 1.150 ;
        RECT 162.650 0.770 163.030 1.150 ;
        RECT 163.310 0.770 163.690 1.150 ;
        RECT 164.230 0.770 164.610 1.150 ;
        RECT 164.890 0.770 165.270 1.150 ;
        RECT 165.550 0.770 165.930 1.150 ;
        RECT 166.310 0.770 166.690 1.150 ;
        RECT 167.630 0.770 168.010 1.150 ;
        RECT 169.830 0.770 170.210 1.150 ;
        RECT 170.490 0.770 170.870 1.150 ;
        RECT 171.150 0.770 171.530 1.150 ;
        RECT 172.070 0.770 172.450 1.150 ;
        RECT 172.730 0.770 173.110 1.150 ;
        RECT 173.390 0.770 173.770 1.150 ;
        RECT 174.410 0.770 174.790 1.150 ;
      LAYER Via2 ;
        RECT 0.815 58.795 1.095 59.075 ;
        RECT 0.815 58.135 1.095 58.415 ;
        RECT 0.815 57.475 1.095 57.755 ;
        RECT 0.815 56.815 1.095 57.095 ;
        RECT 0.815 56.155 1.095 56.435 ;
        RECT 0.815 55.495 1.095 55.775 ;
        RECT 0.815 54.835 1.095 55.115 ;
        RECT 0.815 54.175 1.095 54.455 ;
        RECT 0.815 53.515 1.095 53.795 ;
        RECT 0.815 52.855 1.095 53.135 ;
        RECT 0.815 52.195 1.095 52.475 ;
        RECT 0.815 51.535 1.095 51.815 ;
        RECT 0.815 50.875 1.095 51.155 ;
        RECT 0.815 50.215 1.095 50.495 ;
        RECT 5.300 47.855 5.580 48.135 ;
        RECT 5.960 47.855 6.240 48.135 ;
        RECT 6.620 47.855 6.900 48.135 ;
        RECT 5.300 47.195 5.580 47.475 ;
        RECT 5.960 47.195 6.240 47.475 ;
        RECT 6.620 47.195 6.900 47.475 ;
        RECT 5.300 46.535 5.580 46.815 ;
        RECT 5.960 46.535 6.240 46.815 ;
        RECT 6.620 46.535 6.900 46.815 ;
        RECT 5.300 22.255 5.580 22.535 ;
        RECT 5.960 22.255 6.240 22.535 ;
        RECT 6.620 22.255 6.900 22.535 ;
        RECT 5.300 21.595 5.580 21.875 ;
        RECT 5.960 21.595 6.240 21.875 ;
        RECT 6.620 21.595 6.900 21.875 ;
        RECT 5.300 20.935 5.580 21.215 ;
        RECT 5.960 20.935 6.240 21.215 ;
        RECT 6.620 20.935 6.900 21.215 ;
        RECT 11.105 58.795 11.385 59.075 ;
        RECT 11.105 58.135 11.385 58.415 ;
        RECT 11.105 57.475 11.385 57.755 ;
        RECT 11.105 56.815 11.385 57.095 ;
        RECT 11.105 56.155 11.385 56.435 ;
        RECT 11.105 55.495 11.385 55.775 ;
        RECT 11.105 54.835 11.385 55.115 ;
        RECT 11.105 54.175 11.385 54.455 ;
        RECT 11.105 53.515 11.385 53.795 ;
        RECT 11.105 52.855 11.385 53.135 ;
        RECT 11.105 52.195 11.385 52.475 ;
        RECT 11.105 51.535 11.385 51.815 ;
        RECT 11.105 50.875 11.385 51.155 ;
        RECT 11.105 50.215 11.385 50.495 ;
        RECT 21.390 58.795 21.670 59.075 ;
        RECT 22.810 58.795 23.090 59.075 ;
        RECT 21.390 58.135 21.670 58.415 ;
        RECT 22.810 58.135 23.090 58.415 ;
        RECT 21.390 57.475 21.670 57.755 ;
        RECT 22.810 57.475 23.090 57.755 ;
        RECT 21.390 56.815 21.670 57.095 ;
        RECT 22.810 56.815 23.090 57.095 ;
        RECT 21.390 56.155 21.670 56.435 ;
        RECT 22.810 56.155 23.090 56.435 ;
        RECT 21.390 55.495 21.670 55.775 ;
        RECT 22.810 55.495 23.090 55.775 ;
        RECT 21.390 54.835 21.670 55.115 ;
        RECT 22.810 54.835 23.090 55.115 ;
        RECT 21.390 54.175 21.670 54.455 ;
        RECT 22.810 54.175 23.090 54.455 ;
        RECT 21.390 53.515 21.670 53.795 ;
        RECT 22.810 53.515 23.090 53.795 ;
        RECT 21.390 52.855 21.670 53.135 ;
        RECT 22.810 52.855 23.090 53.135 ;
        RECT 21.390 52.195 21.670 52.475 ;
        RECT 22.810 52.195 23.090 52.475 ;
        RECT 21.390 51.535 21.670 51.815 ;
        RECT 22.810 51.535 23.090 51.815 ;
        RECT 21.390 50.875 21.670 51.155 ;
        RECT 22.810 50.875 23.090 51.155 ;
        RECT 21.390 50.215 21.670 50.495 ;
        RECT 22.810 50.215 23.090 50.495 ;
        RECT 27.295 47.855 27.575 48.135 ;
        RECT 27.955 47.855 28.235 48.135 ;
        RECT 28.615 47.855 28.895 48.135 ;
        RECT 27.295 47.195 27.575 47.475 ;
        RECT 27.955 47.195 28.235 47.475 ;
        RECT 28.615 47.195 28.895 47.475 ;
        RECT 27.295 46.535 27.575 46.815 ;
        RECT 27.955 46.535 28.235 46.815 ;
        RECT 28.615 46.535 28.895 46.815 ;
        RECT 15.600 45.155 15.880 45.435 ;
        RECT 16.260 45.155 16.540 45.435 ;
        RECT 16.920 45.155 17.200 45.435 ;
        RECT 15.600 44.495 15.880 44.775 ;
        RECT 16.260 44.495 16.540 44.775 ;
        RECT 16.920 44.495 17.200 44.775 ;
        RECT 15.600 43.835 15.880 44.115 ;
        RECT 16.260 43.835 16.540 44.115 ;
        RECT 16.920 43.835 17.200 44.115 ;
        RECT 15.600 24.955 15.880 25.235 ;
        RECT 16.260 24.955 16.540 25.235 ;
        RECT 16.920 24.955 17.200 25.235 ;
        RECT 15.600 24.295 15.880 24.575 ;
        RECT 16.260 24.295 16.540 24.575 ;
        RECT 16.920 24.295 17.200 24.575 ;
        RECT 15.600 23.635 15.880 23.915 ;
        RECT 16.260 23.635 16.540 23.915 ;
        RECT 16.920 23.635 17.200 23.915 ;
        RECT 27.295 22.255 27.575 22.535 ;
        RECT 27.955 22.255 28.235 22.535 ;
        RECT 28.615 22.255 28.895 22.535 ;
        RECT 27.295 21.595 27.575 21.875 ;
        RECT 27.955 21.595 28.235 21.875 ;
        RECT 28.615 21.595 28.895 21.875 ;
        RECT 27.295 20.935 27.575 21.215 ;
        RECT 27.955 20.935 28.235 21.215 ;
        RECT 28.615 20.935 28.895 21.215 ;
        RECT 33.100 58.795 33.380 59.075 ;
        RECT 33.100 58.135 33.380 58.415 ;
        RECT 33.100 57.475 33.380 57.755 ;
        RECT 33.100 56.815 33.380 57.095 ;
        RECT 33.100 56.155 33.380 56.435 ;
        RECT 33.100 55.495 33.380 55.775 ;
        RECT 33.100 54.835 33.380 55.115 ;
        RECT 33.100 54.175 33.380 54.455 ;
        RECT 33.100 53.515 33.380 53.795 ;
        RECT 33.100 52.855 33.380 53.135 ;
        RECT 33.100 52.195 33.380 52.475 ;
        RECT 33.100 51.535 33.380 51.815 ;
        RECT 33.100 50.875 33.380 51.155 ;
        RECT 33.100 50.215 33.380 50.495 ;
        RECT 43.385 58.795 43.665 59.075 ;
        RECT 44.805 58.795 45.085 59.075 ;
        RECT 43.385 58.135 43.665 58.415 ;
        RECT 44.805 58.135 45.085 58.415 ;
        RECT 43.385 57.475 43.665 57.755 ;
        RECT 44.805 57.475 45.085 57.755 ;
        RECT 43.385 56.815 43.665 57.095 ;
        RECT 44.805 56.815 45.085 57.095 ;
        RECT 43.385 56.155 43.665 56.435 ;
        RECT 44.805 56.155 45.085 56.435 ;
        RECT 43.385 55.495 43.665 55.775 ;
        RECT 44.805 55.495 45.085 55.775 ;
        RECT 43.385 54.835 43.665 55.115 ;
        RECT 44.805 54.835 45.085 55.115 ;
        RECT 43.385 54.175 43.665 54.455 ;
        RECT 44.805 54.175 45.085 54.455 ;
        RECT 43.385 53.515 43.665 53.795 ;
        RECT 44.805 53.515 45.085 53.795 ;
        RECT 43.385 52.855 43.665 53.135 ;
        RECT 44.805 52.855 45.085 53.135 ;
        RECT 43.385 52.195 43.665 52.475 ;
        RECT 44.805 52.195 45.085 52.475 ;
        RECT 43.385 51.535 43.665 51.815 ;
        RECT 44.805 51.535 45.085 51.815 ;
        RECT 43.385 50.875 43.665 51.155 ;
        RECT 44.805 50.875 45.085 51.155 ;
        RECT 43.385 50.215 43.665 50.495 ;
        RECT 44.805 50.215 45.085 50.495 ;
        RECT 49.290 47.855 49.570 48.135 ;
        RECT 49.950 47.855 50.230 48.135 ;
        RECT 50.610 47.855 50.890 48.135 ;
        RECT 49.290 47.195 49.570 47.475 ;
        RECT 49.950 47.195 50.230 47.475 ;
        RECT 50.610 47.195 50.890 47.475 ;
        RECT 49.290 46.535 49.570 46.815 ;
        RECT 49.950 46.535 50.230 46.815 ;
        RECT 50.610 46.535 50.890 46.815 ;
        RECT 37.595 45.155 37.875 45.435 ;
        RECT 38.255 45.155 38.535 45.435 ;
        RECT 38.915 45.155 39.195 45.435 ;
        RECT 37.595 44.495 37.875 44.775 ;
        RECT 38.255 44.495 38.535 44.775 ;
        RECT 38.915 44.495 39.195 44.775 ;
        RECT 37.595 43.835 37.875 44.115 ;
        RECT 38.255 43.835 38.535 44.115 ;
        RECT 38.915 43.835 39.195 44.115 ;
        RECT 37.595 24.955 37.875 25.235 ;
        RECT 38.255 24.955 38.535 25.235 ;
        RECT 38.915 24.955 39.195 25.235 ;
        RECT 37.595 24.295 37.875 24.575 ;
        RECT 38.255 24.295 38.535 24.575 ;
        RECT 38.915 24.295 39.195 24.575 ;
        RECT 37.595 23.635 37.875 23.915 ;
        RECT 38.255 23.635 38.535 23.915 ;
        RECT 38.915 23.635 39.195 23.915 ;
        RECT 49.290 22.255 49.570 22.535 ;
        RECT 49.950 22.255 50.230 22.535 ;
        RECT 50.610 22.255 50.890 22.535 ;
        RECT 49.290 21.595 49.570 21.875 ;
        RECT 49.950 21.595 50.230 21.875 ;
        RECT 50.610 21.595 50.890 21.875 ;
        RECT 49.290 20.935 49.570 21.215 ;
        RECT 49.950 20.935 50.230 21.215 ;
        RECT 50.610 20.935 50.890 21.215 ;
        RECT 55.095 58.795 55.375 59.075 ;
        RECT 55.095 58.135 55.375 58.415 ;
        RECT 55.095 57.475 55.375 57.755 ;
        RECT 55.095 56.815 55.375 57.095 ;
        RECT 55.095 56.155 55.375 56.435 ;
        RECT 55.095 55.495 55.375 55.775 ;
        RECT 55.095 54.835 55.375 55.115 ;
        RECT 55.095 54.175 55.375 54.455 ;
        RECT 55.095 53.515 55.375 53.795 ;
        RECT 55.095 52.855 55.375 53.135 ;
        RECT 55.095 52.195 55.375 52.475 ;
        RECT 55.095 51.535 55.375 51.815 ;
        RECT 55.095 50.875 55.375 51.155 ;
        RECT 55.095 50.215 55.375 50.495 ;
        RECT 65.380 58.795 65.660 59.075 ;
        RECT 66.800 58.795 67.080 59.075 ;
        RECT 65.380 58.135 65.660 58.415 ;
        RECT 66.800 58.135 67.080 58.415 ;
        RECT 65.380 57.475 65.660 57.755 ;
        RECT 66.800 57.475 67.080 57.755 ;
        RECT 65.380 56.815 65.660 57.095 ;
        RECT 66.800 56.815 67.080 57.095 ;
        RECT 65.380 56.155 65.660 56.435 ;
        RECT 66.800 56.155 67.080 56.435 ;
        RECT 65.380 55.495 65.660 55.775 ;
        RECT 66.800 55.495 67.080 55.775 ;
        RECT 65.380 54.835 65.660 55.115 ;
        RECT 66.800 54.835 67.080 55.115 ;
        RECT 65.380 54.175 65.660 54.455 ;
        RECT 66.800 54.175 67.080 54.455 ;
        RECT 65.380 53.515 65.660 53.795 ;
        RECT 66.800 53.515 67.080 53.795 ;
        RECT 65.380 52.855 65.660 53.135 ;
        RECT 66.800 52.855 67.080 53.135 ;
        RECT 65.380 52.195 65.660 52.475 ;
        RECT 66.800 52.195 67.080 52.475 ;
        RECT 65.380 51.535 65.660 51.815 ;
        RECT 66.800 51.535 67.080 51.815 ;
        RECT 65.380 50.875 65.660 51.155 ;
        RECT 66.800 50.875 67.080 51.155 ;
        RECT 65.380 50.215 65.660 50.495 ;
        RECT 66.800 50.215 67.080 50.495 ;
        RECT 71.285 47.855 71.565 48.135 ;
        RECT 71.945 47.855 72.225 48.135 ;
        RECT 72.605 47.855 72.885 48.135 ;
        RECT 71.285 47.195 71.565 47.475 ;
        RECT 71.945 47.195 72.225 47.475 ;
        RECT 72.605 47.195 72.885 47.475 ;
        RECT 71.285 46.535 71.565 46.815 ;
        RECT 71.945 46.535 72.225 46.815 ;
        RECT 72.605 46.535 72.885 46.815 ;
        RECT 59.590 45.155 59.870 45.435 ;
        RECT 60.250 45.155 60.530 45.435 ;
        RECT 60.910 45.155 61.190 45.435 ;
        RECT 59.590 44.495 59.870 44.775 ;
        RECT 60.250 44.495 60.530 44.775 ;
        RECT 60.910 44.495 61.190 44.775 ;
        RECT 59.590 43.835 59.870 44.115 ;
        RECT 60.250 43.835 60.530 44.115 ;
        RECT 60.910 43.835 61.190 44.115 ;
        RECT 59.590 24.955 59.870 25.235 ;
        RECT 60.250 24.955 60.530 25.235 ;
        RECT 60.910 24.955 61.190 25.235 ;
        RECT 59.590 24.295 59.870 24.575 ;
        RECT 60.250 24.295 60.530 24.575 ;
        RECT 60.910 24.295 61.190 24.575 ;
        RECT 59.590 23.635 59.870 23.915 ;
        RECT 60.250 23.635 60.530 23.915 ;
        RECT 60.910 23.635 61.190 23.915 ;
        RECT 71.285 22.255 71.565 22.535 ;
        RECT 71.945 22.255 72.225 22.535 ;
        RECT 72.605 22.255 72.885 22.535 ;
        RECT 71.285 21.595 71.565 21.875 ;
        RECT 71.945 21.595 72.225 21.875 ;
        RECT 72.605 21.595 72.885 21.875 ;
        RECT 71.285 20.935 71.565 21.215 ;
        RECT 71.945 20.935 72.225 21.215 ;
        RECT 72.605 20.935 72.885 21.215 ;
        RECT 77.090 58.795 77.370 59.075 ;
        RECT 77.090 58.135 77.370 58.415 ;
        RECT 77.090 57.475 77.370 57.755 ;
        RECT 77.090 56.815 77.370 57.095 ;
        RECT 77.090 56.155 77.370 56.435 ;
        RECT 77.090 55.495 77.370 55.775 ;
        RECT 77.090 54.835 77.370 55.115 ;
        RECT 77.090 54.175 77.370 54.455 ;
        RECT 77.090 53.515 77.370 53.795 ;
        RECT 77.090 52.855 77.370 53.135 ;
        RECT 77.090 52.195 77.370 52.475 ;
        RECT 77.090 51.535 77.370 51.815 ;
        RECT 77.090 50.875 77.370 51.155 ;
        RECT 77.090 50.215 77.370 50.495 ;
        RECT 87.375 58.795 87.655 59.075 ;
        RECT 88.795 58.795 89.075 59.075 ;
        RECT 87.375 58.135 87.655 58.415 ;
        RECT 88.795 58.135 89.075 58.415 ;
        RECT 87.375 57.475 87.655 57.755 ;
        RECT 88.795 57.475 89.075 57.755 ;
        RECT 87.375 56.815 87.655 57.095 ;
        RECT 88.795 56.815 89.075 57.095 ;
        RECT 87.375 56.155 87.655 56.435 ;
        RECT 88.795 56.155 89.075 56.435 ;
        RECT 87.375 55.495 87.655 55.775 ;
        RECT 88.795 55.495 89.075 55.775 ;
        RECT 87.375 54.835 87.655 55.115 ;
        RECT 88.795 54.835 89.075 55.115 ;
        RECT 87.375 54.175 87.655 54.455 ;
        RECT 88.795 54.175 89.075 54.455 ;
        RECT 87.375 53.515 87.655 53.795 ;
        RECT 88.795 53.515 89.075 53.795 ;
        RECT 87.375 52.855 87.655 53.135 ;
        RECT 88.795 52.855 89.075 53.135 ;
        RECT 87.375 52.195 87.655 52.475 ;
        RECT 88.795 52.195 89.075 52.475 ;
        RECT 87.375 51.535 87.655 51.815 ;
        RECT 88.795 51.535 89.075 51.815 ;
        RECT 87.375 50.875 87.655 51.155 ;
        RECT 88.795 50.875 89.075 51.155 ;
        RECT 87.375 50.215 87.655 50.495 ;
        RECT 88.795 50.215 89.075 50.495 ;
        RECT 93.280 47.855 93.560 48.135 ;
        RECT 93.940 47.855 94.220 48.135 ;
        RECT 94.600 47.855 94.880 48.135 ;
        RECT 93.280 47.195 93.560 47.475 ;
        RECT 93.940 47.195 94.220 47.475 ;
        RECT 94.600 47.195 94.880 47.475 ;
        RECT 93.280 46.535 93.560 46.815 ;
        RECT 93.940 46.535 94.220 46.815 ;
        RECT 94.600 46.535 94.880 46.815 ;
        RECT 81.585 45.155 81.865 45.435 ;
        RECT 82.245 45.155 82.525 45.435 ;
        RECT 82.905 45.155 83.185 45.435 ;
        RECT 81.585 44.495 81.865 44.775 ;
        RECT 82.245 44.495 82.525 44.775 ;
        RECT 82.905 44.495 83.185 44.775 ;
        RECT 81.585 43.835 81.865 44.115 ;
        RECT 82.245 43.835 82.525 44.115 ;
        RECT 82.905 43.835 83.185 44.115 ;
        RECT 81.585 24.955 81.865 25.235 ;
        RECT 82.245 24.955 82.525 25.235 ;
        RECT 82.905 24.955 83.185 25.235 ;
        RECT 81.585 24.295 81.865 24.575 ;
        RECT 82.245 24.295 82.525 24.575 ;
        RECT 82.905 24.295 83.185 24.575 ;
        RECT 81.585 23.635 81.865 23.915 ;
        RECT 82.245 23.635 82.525 23.915 ;
        RECT 82.905 23.635 83.185 23.915 ;
        RECT 93.280 22.255 93.560 22.535 ;
        RECT 93.940 22.255 94.220 22.535 ;
        RECT 94.600 22.255 94.880 22.535 ;
        RECT 93.280 21.595 93.560 21.875 ;
        RECT 93.940 21.595 94.220 21.875 ;
        RECT 94.600 21.595 94.880 21.875 ;
        RECT 93.280 20.935 93.560 21.215 ;
        RECT 93.940 20.935 94.220 21.215 ;
        RECT 94.600 20.935 94.880 21.215 ;
        RECT 99.085 58.795 99.365 59.075 ;
        RECT 99.085 58.135 99.365 58.415 ;
        RECT 99.085 57.475 99.365 57.755 ;
        RECT 99.085 56.815 99.365 57.095 ;
        RECT 99.085 56.155 99.365 56.435 ;
        RECT 99.085 55.495 99.365 55.775 ;
        RECT 99.085 54.835 99.365 55.115 ;
        RECT 99.085 54.175 99.365 54.455 ;
        RECT 99.085 53.515 99.365 53.795 ;
        RECT 99.085 52.855 99.365 53.135 ;
        RECT 99.085 52.195 99.365 52.475 ;
        RECT 99.085 51.535 99.365 51.815 ;
        RECT 99.085 50.875 99.365 51.155 ;
        RECT 99.085 50.215 99.365 50.495 ;
        RECT 109.370 58.795 109.650 59.075 ;
        RECT 110.790 58.795 111.070 59.075 ;
        RECT 109.370 58.135 109.650 58.415 ;
        RECT 110.790 58.135 111.070 58.415 ;
        RECT 109.370 57.475 109.650 57.755 ;
        RECT 110.790 57.475 111.070 57.755 ;
        RECT 109.370 56.815 109.650 57.095 ;
        RECT 110.790 56.815 111.070 57.095 ;
        RECT 109.370 56.155 109.650 56.435 ;
        RECT 110.790 56.155 111.070 56.435 ;
        RECT 109.370 55.495 109.650 55.775 ;
        RECT 110.790 55.495 111.070 55.775 ;
        RECT 109.370 54.835 109.650 55.115 ;
        RECT 110.790 54.835 111.070 55.115 ;
        RECT 109.370 54.175 109.650 54.455 ;
        RECT 110.790 54.175 111.070 54.455 ;
        RECT 109.370 53.515 109.650 53.795 ;
        RECT 110.790 53.515 111.070 53.795 ;
        RECT 109.370 52.855 109.650 53.135 ;
        RECT 110.790 52.855 111.070 53.135 ;
        RECT 109.370 52.195 109.650 52.475 ;
        RECT 110.790 52.195 111.070 52.475 ;
        RECT 109.370 51.535 109.650 51.815 ;
        RECT 110.790 51.535 111.070 51.815 ;
        RECT 109.370 50.875 109.650 51.155 ;
        RECT 110.790 50.875 111.070 51.155 ;
        RECT 109.370 50.215 109.650 50.495 ;
        RECT 110.790 50.215 111.070 50.495 ;
        RECT 115.275 47.855 115.555 48.135 ;
        RECT 115.935 47.855 116.215 48.135 ;
        RECT 116.595 47.855 116.875 48.135 ;
        RECT 115.275 47.195 115.555 47.475 ;
        RECT 115.935 47.195 116.215 47.475 ;
        RECT 116.595 47.195 116.875 47.475 ;
        RECT 115.275 46.535 115.555 46.815 ;
        RECT 115.935 46.535 116.215 46.815 ;
        RECT 116.595 46.535 116.875 46.815 ;
        RECT 103.580 45.155 103.860 45.435 ;
        RECT 104.240 45.155 104.520 45.435 ;
        RECT 104.900 45.155 105.180 45.435 ;
        RECT 103.580 44.495 103.860 44.775 ;
        RECT 104.240 44.495 104.520 44.775 ;
        RECT 104.900 44.495 105.180 44.775 ;
        RECT 103.580 43.835 103.860 44.115 ;
        RECT 104.240 43.835 104.520 44.115 ;
        RECT 104.900 43.835 105.180 44.115 ;
        RECT 103.580 24.955 103.860 25.235 ;
        RECT 104.240 24.955 104.520 25.235 ;
        RECT 104.900 24.955 105.180 25.235 ;
        RECT 103.580 24.295 103.860 24.575 ;
        RECT 104.240 24.295 104.520 24.575 ;
        RECT 104.900 24.295 105.180 24.575 ;
        RECT 103.580 23.635 103.860 23.915 ;
        RECT 104.240 23.635 104.520 23.915 ;
        RECT 104.900 23.635 105.180 23.915 ;
        RECT 115.275 22.255 115.555 22.535 ;
        RECT 115.935 22.255 116.215 22.535 ;
        RECT 116.595 22.255 116.875 22.535 ;
        RECT 115.275 21.595 115.555 21.875 ;
        RECT 115.935 21.595 116.215 21.875 ;
        RECT 116.595 21.595 116.875 21.875 ;
        RECT 115.275 20.935 115.555 21.215 ;
        RECT 115.935 20.935 116.215 21.215 ;
        RECT 116.595 20.935 116.875 21.215 ;
        RECT 121.080 58.795 121.360 59.075 ;
        RECT 121.080 58.135 121.360 58.415 ;
        RECT 121.080 57.475 121.360 57.755 ;
        RECT 121.080 56.815 121.360 57.095 ;
        RECT 121.080 56.155 121.360 56.435 ;
        RECT 121.080 55.495 121.360 55.775 ;
        RECT 121.080 54.835 121.360 55.115 ;
        RECT 121.080 54.175 121.360 54.455 ;
        RECT 121.080 53.515 121.360 53.795 ;
        RECT 121.080 52.855 121.360 53.135 ;
        RECT 121.080 52.195 121.360 52.475 ;
        RECT 121.080 51.535 121.360 51.815 ;
        RECT 121.080 50.875 121.360 51.155 ;
        RECT 121.080 50.215 121.360 50.495 ;
        RECT 131.365 58.795 131.645 59.075 ;
        RECT 132.785 58.795 133.065 59.075 ;
        RECT 131.365 58.135 131.645 58.415 ;
        RECT 132.785 58.135 133.065 58.415 ;
        RECT 131.365 57.475 131.645 57.755 ;
        RECT 132.785 57.475 133.065 57.755 ;
        RECT 131.365 56.815 131.645 57.095 ;
        RECT 132.785 56.815 133.065 57.095 ;
        RECT 131.365 56.155 131.645 56.435 ;
        RECT 132.785 56.155 133.065 56.435 ;
        RECT 131.365 55.495 131.645 55.775 ;
        RECT 132.785 55.495 133.065 55.775 ;
        RECT 131.365 54.835 131.645 55.115 ;
        RECT 132.785 54.835 133.065 55.115 ;
        RECT 131.365 54.175 131.645 54.455 ;
        RECT 132.785 54.175 133.065 54.455 ;
        RECT 131.365 53.515 131.645 53.795 ;
        RECT 132.785 53.515 133.065 53.795 ;
        RECT 131.365 52.855 131.645 53.135 ;
        RECT 132.785 52.855 133.065 53.135 ;
        RECT 131.365 52.195 131.645 52.475 ;
        RECT 132.785 52.195 133.065 52.475 ;
        RECT 131.365 51.535 131.645 51.815 ;
        RECT 132.785 51.535 133.065 51.815 ;
        RECT 131.365 50.875 131.645 51.155 ;
        RECT 132.785 50.875 133.065 51.155 ;
        RECT 131.365 50.215 131.645 50.495 ;
        RECT 132.785 50.215 133.065 50.495 ;
        RECT 137.270 47.855 137.550 48.135 ;
        RECT 137.930 47.855 138.210 48.135 ;
        RECT 138.590 47.855 138.870 48.135 ;
        RECT 137.270 47.195 137.550 47.475 ;
        RECT 137.930 47.195 138.210 47.475 ;
        RECT 138.590 47.195 138.870 47.475 ;
        RECT 137.270 46.535 137.550 46.815 ;
        RECT 137.930 46.535 138.210 46.815 ;
        RECT 138.590 46.535 138.870 46.815 ;
        RECT 125.575 45.155 125.855 45.435 ;
        RECT 126.235 45.155 126.515 45.435 ;
        RECT 126.895 45.155 127.175 45.435 ;
        RECT 125.575 44.495 125.855 44.775 ;
        RECT 126.235 44.495 126.515 44.775 ;
        RECT 126.895 44.495 127.175 44.775 ;
        RECT 125.575 43.835 125.855 44.115 ;
        RECT 126.235 43.835 126.515 44.115 ;
        RECT 126.895 43.835 127.175 44.115 ;
        RECT 125.575 24.955 125.855 25.235 ;
        RECT 126.235 24.955 126.515 25.235 ;
        RECT 126.895 24.955 127.175 25.235 ;
        RECT 125.575 24.295 125.855 24.575 ;
        RECT 126.235 24.295 126.515 24.575 ;
        RECT 126.895 24.295 127.175 24.575 ;
        RECT 125.575 23.635 125.855 23.915 ;
        RECT 126.235 23.635 126.515 23.915 ;
        RECT 126.895 23.635 127.175 23.915 ;
        RECT 137.270 22.255 137.550 22.535 ;
        RECT 137.930 22.255 138.210 22.535 ;
        RECT 138.590 22.255 138.870 22.535 ;
        RECT 137.270 21.595 137.550 21.875 ;
        RECT 137.930 21.595 138.210 21.875 ;
        RECT 138.590 21.595 138.870 21.875 ;
        RECT 137.270 20.935 137.550 21.215 ;
        RECT 137.930 20.935 138.210 21.215 ;
        RECT 138.590 20.935 138.870 21.215 ;
        RECT 143.075 58.795 143.355 59.075 ;
        RECT 143.075 58.135 143.355 58.415 ;
        RECT 143.075 57.475 143.355 57.755 ;
        RECT 143.075 56.815 143.355 57.095 ;
        RECT 143.075 56.155 143.355 56.435 ;
        RECT 143.075 55.495 143.355 55.775 ;
        RECT 143.075 54.835 143.355 55.115 ;
        RECT 143.075 54.175 143.355 54.455 ;
        RECT 143.075 53.515 143.355 53.795 ;
        RECT 143.075 52.855 143.355 53.135 ;
        RECT 143.075 52.195 143.355 52.475 ;
        RECT 143.075 51.535 143.355 51.815 ;
        RECT 143.075 50.875 143.355 51.155 ;
        RECT 143.075 50.215 143.355 50.495 ;
        RECT 153.360 58.795 153.640 59.075 ;
        RECT 154.780 58.795 155.060 59.075 ;
        RECT 153.360 58.135 153.640 58.415 ;
        RECT 154.780 58.135 155.060 58.415 ;
        RECT 153.360 57.475 153.640 57.755 ;
        RECT 154.780 57.475 155.060 57.755 ;
        RECT 153.360 56.815 153.640 57.095 ;
        RECT 154.780 56.815 155.060 57.095 ;
        RECT 153.360 56.155 153.640 56.435 ;
        RECT 154.780 56.155 155.060 56.435 ;
        RECT 153.360 55.495 153.640 55.775 ;
        RECT 154.780 55.495 155.060 55.775 ;
        RECT 153.360 54.835 153.640 55.115 ;
        RECT 154.780 54.835 155.060 55.115 ;
        RECT 153.360 54.175 153.640 54.455 ;
        RECT 154.780 54.175 155.060 54.455 ;
        RECT 153.360 53.515 153.640 53.795 ;
        RECT 154.780 53.515 155.060 53.795 ;
        RECT 153.360 52.855 153.640 53.135 ;
        RECT 154.780 52.855 155.060 53.135 ;
        RECT 153.360 52.195 153.640 52.475 ;
        RECT 154.780 52.195 155.060 52.475 ;
        RECT 153.360 51.535 153.640 51.815 ;
        RECT 154.780 51.535 155.060 51.815 ;
        RECT 153.360 50.875 153.640 51.155 ;
        RECT 154.780 50.875 155.060 51.155 ;
        RECT 153.360 50.215 153.640 50.495 ;
        RECT 154.780 50.215 155.060 50.495 ;
        RECT 159.265 47.855 159.545 48.135 ;
        RECT 159.925 47.855 160.205 48.135 ;
        RECT 160.585 47.855 160.865 48.135 ;
        RECT 159.265 47.195 159.545 47.475 ;
        RECT 159.925 47.195 160.205 47.475 ;
        RECT 160.585 47.195 160.865 47.475 ;
        RECT 159.265 46.535 159.545 46.815 ;
        RECT 159.925 46.535 160.205 46.815 ;
        RECT 160.585 46.535 160.865 46.815 ;
        RECT 147.570 45.155 147.850 45.435 ;
        RECT 148.230 45.155 148.510 45.435 ;
        RECT 148.890 45.155 149.170 45.435 ;
        RECT 147.570 44.495 147.850 44.775 ;
        RECT 148.230 44.495 148.510 44.775 ;
        RECT 148.890 44.495 149.170 44.775 ;
        RECT 147.570 43.835 147.850 44.115 ;
        RECT 148.230 43.835 148.510 44.115 ;
        RECT 148.890 43.835 149.170 44.115 ;
        RECT 147.570 24.955 147.850 25.235 ;
        RECT 148.230 24.955 148.510 25.235 ;
        RECT 148.890 24.955 149.170 25.235 ;
        RECT 147.570 24.295 147.850 24.575 ;
        RECT 148.230 24.295 148.510 24.575 ;
        RECT 148.890 24.295 149.170 24.575 ;
        RECT 147.570 23.635 147.850 23.915 ;
        RECT 148.230 23.635 148.510 23.915 ;
        RECT 148.890 23.635 149.170 23.915 ;
        RECT 159.265 22.255 159.545 22.535 ;
        RECT 159.925 22.255 160.205 22.535 ;
        RECT 160.585 22.255 160.865 22.535 ;
        RECT 159.265 21.595 159.545 21.875 ;
        RECT 159.925 21.595 160.205 21.875 ;
        RECT 160.585 21.595 160.865 21.875 ;
        RECT 159.265 20.935 159.545 21.215 ;
        RECT 159.925 20.935 160.205 21.215 ;
        RECT 160.585 20.935 160.865 21.215 ;
        RECT 165.070 58.795 165.350 59.075 ;
        RECT 165.070 58.135 165.350 58.415 ;
        RECT 165.070 57.475 165.350 57.755 ;
        RECT 165.070 56.815 165.350 57.095 ;
        RECT 165.070 56.155 165.350 56.435 ;
        RECT 165.070 55.495 165.350 55.775 ;
        RECT 165.070 54.835 165.350 55.115 ;
        RECT 165.070 54.175 165.350 54.455 ;
        RECT 165.070 53.515 165.350 53.795 ;
        RECT 165.070 52.855 165.350 53.135 ;
        RECT 165.070 52.195 165.350 52.475 ;
        RECT 165.070 51.535 165.350 51.815 ;
        RECT 165.070 50.875 165.350 51.155 ;
        RECT 165.070 50.215 165.350 50.495 ;
        RECT 175.355 58.795 175.635 59.075 ;
        RECT 175.355 58.135 175.635 58.415 ;
        RECT 175.355 57.475 175.635 57.755 ;
        RECT 175.355 56.815 175.635 57.095 ;
        RECT 175.355 56.155 175.635 56.435 ;
        RECT 175.355 55.495 175.635 55.775 ;
        RECT 177.200 55.165 177.480 55.445 ;
        RECT 178.985 55.165 179.265 55.445 ;
        RECT 181.840 55.165 182.120 55.445 ;
        RECT 183.625 55.165 183.905 55.445 ;
        RECT 186.480 55.165 186.760 55.445 ;
        RECT 188.265 55.165 188.545 55.445 ;
        RECT 191.120 55.165 191.400 55.445 ;
        RECT 192.905 55.165 193.185 55.445 ;
        RECT 175.355 54.835 175.635 55.115 ;
        RECT 177.200 54.505 177.480 54.785 ;
        RECT 178.985 54.505 179.265 54.785 ;
        RECT 181.840 54.505 182.120 54.785 ;
        RECT 183.625 54.505 183.905 54.785 ;
        RECT 186.480 54.505 186.760 54.785 ;
        RECT 188.265 54.505 188.545 54.785 ;
        RECT 191.120 54.505 191.400 54.785 ;
        RECT 192.905 54.505 193.185 54.785 ;
        RECT 175.355 54.175 175.635 54.455 ;
        RECT 177.200 53.845 177.480 54.125 ;
        RECT 178.985 53.845 179.265 54.125 ;
        RECT 181.840 53.845 182.120 54.125 ;
        RECT 183.625 53.845 183.905 54.125 ;
        RECT 186.480 53.845 186.760 54.125 ;
        RECT 188.265 53.845 188.545 54.125 ;
        RECT 191.120 53.845 191.400 54.125 ;
        RECT 192.905 53.845 193.185 54.125 ;
        RECT 175.355 53.515 175.635 53.795 ;
        RECT 177.200 53.185 177.480 53.465 ;
        RECT 178.985 53.185 179.265 53.465 ;
        RECT 181.840 53.185 182.120 53.465 ;
        RECT 183.625 53.185 183.905 53.465 ;
        RECT 186.480 53.185 186.760 53.465 ;
        RECT 188.265 53.185 188.545 53.465 ;
        RECT 191.120 53.185 191.400 53.465 ;
        RECT 192.905 53.185 193.185 53.465 ;
        RECT 175.355 52.855 175.635 53.135 ;
        RECT 177.200 52.525 177.480 52.805 ;
        RECT 178.985 52.525 179.265 52.805 ;
        RECT 181.840 52.525 182.120 52.805 ;
        RECT 183.625 52.525 183.905 52.805 ;
        RECT 186.480 52.525 186.760 52.805 ;
        RECT 188.265 52.525 188.545 52.805 ;
        RECT 191.120 52.525 191.400 52.805 ;
        RECT 192.905 52.525 193.185 52.805 ;
        RECT 175.355 52.195 175.635 52.475 ;
        RECT 177.200 51.865 177.480 52.145 ;
        RECT 178.985 51.865 179.265 52.145 ;
        RECT 181.840 51.865 182.120 52.145 ;
        RECT 183.625 51.865 183.905 52.145 ;
        RECT 186.480 51.865 186.760 52.145 ;
        RECT 188.265 51.865 188.545 52.145 ;
        RECT 191.120 51.865 191.400 52.145 ;
        RECT 192.905 51.865 193.185 52.145 ;
        RECT 175.355 51.535 175.635 51.815 ;
        RECT 177.200 51.205 177.480 51.485 ;
        RECT 178.985 51.205 179.265 51.485 ;
        RECT 181.840 51.205 182.120 51.485 ;
        RECT 183.625 51.205 183.905 51.485 ;
        RECT 186.480 51.205 186.760 51.485 ;
        RECT 188.265 51.205 188.545 51.485 ;
        RECT 191.120 51.205 191.400 51.485 ;
        RECT 192.905 51.205 193.185 51.485 ;
        RECT 175.355 50.875 175.635 51.155 ;
        RECT 177.200 50.545 177.480 50.825 ;
        RECT 178.985 50.545 179.265 50.825 ;
        RECT 181.840 50.545 182.120 50.825 ;
        RECT 183.625 50.545 183.905 50.825 ;
        RECT 186.480 50.545 186.760 50.825 ;
        RECT 188.265 50.545 188.545 50.825 ;
        RECT 191.120 50.545 191.400 50.825 ;
        RECT 192.905 50.545 193.185 50.825 ;
        RECT 175.355 50.215 175.635 50.495 ;
        RECT 177.960 47.855 178.240 48.135 ;
        RECT 177.960 47.195 178.240 47.475 ;
        RECT 177.960 46.535 178.240 46.815 ;
        RECT 169.565 45.155 169.845 45.435 ;
        RECT 170.225 45.155 170.505 45.435 ;
        RECT 170.885 45.155 171.165 45.435 ;
        RECT 191.880 45.155 192.160 45.435 ;
        RECT 169.565 44.495 169.845 44.775 ;
        RECT 170.225 44.495 170.505 44.775 ;
        RECT 170.885 44.495 171.165 44.775 ;
        RECT 191.880 44.495 192.160 44.775 ;
        RECT 169.565 43.835 169.845 44.115 ;
        RECT 170.225 43.835 170.505 44.115 ;
        RECT 170.885 43.835 171.165 44.115 ;
        RECT 191.880 43.835 192.160 44.115 ;
        RECT 169.565 24.955 169.845 25.235 ;
        RECT 170.225 24.955 170.505 25.235 ;
        RECT 170.885 24.955 171.165 25.235 ;
        RECT 187.240 24.955 187.520 25.235 ;
        RECT 169.565 24.295 169.845 24.575 ;
        RECT 170.225 24.295 170.505 24.575 ;
        RECT 170.885 24.295 171.165 24.575 ;
        RECT 187.240 24.295 187.520 24.575 ;
        RECT 169.565 23.635 169.845 23.915 ;
        RECT 170.225 23.635 170.505 23.915 ;
        RECT 170.885 23.635 171.165 23.915 ;
        RECT 187.240 23.635 187.520 23.915 ;
        RECT 182.600 22.255 182.880 22.535 ;
        RECT 182.600 21.595 182.880 21.875 ;
        RECT 182.600 20.935 182.880 21.215 ;
        RECT 177.200 18.165 177.480 18.445 ;
        RECT 178.985 18.165 179.265 18.445 ;
        RECT 181.840 18.165 182.120 18.445 ;
        RECT 183.625 18.165 183.905 18.445 ;
        RECT 186.480 18.165 186.760 18.445 ;
        RECT 188.265 18.165 188.545 18.445 ;
        RECT 191.120 18.165 191.400 18.445 ;
        RECT 192.905 18.165 193.185 18.445 ;
        RECT 177.200 17.505 177.480 17.785 ;
        RECT 178.985 17.505 179.265 17.785 ;
        RECT 181.840 17.505 182.120 17.785 ;
        RECT 183.625 17.505 183.905 17.785 ;
        RECT 186.480 17.505 186.760 17.785 ;
        RECT 188.265 17.505 188.545 17.785 ;
        RECT 191.120 17.505 191.400 17.785 ;
        RECT 192.905 17.505 193.185 17.785 ;
        RECT 177.200 16.845 177.480 17.125 ;
        RECT 178.985 16.845 179.265 17.125 ;
        RECT 181.840 16.845 182.120 17.125 ;
        RECT 183.625 16.845 183.905 17.125 ;
        RECT 186.480 16.845 186.760 17.125 ;
        RECT 188.265 16.845 188.545 17.125 ;
        RECT 191.120 16.845 191.400 17.125 ;
        RECT 192.905 16.845 193.185 17.125 ;
        RECT 177.200 16.185 177.480 16.465 ;
        RECT 178.985 16.185 179.265 16.465 ;
        RECT 181.840 16.185 182.120 16.465 ;
        RECT 183.625 16.185 183.905 16.465 ;
        RECT 186.480 16.185 186.760 16.465 ;
        RECT 188.265 16.185 188.545 16.465 ;
        RECT 191.120 16.185 191.400 16.465 ;
        RECT 192.905 16.185 193.185 16.465 ;
        RECT 177.200 15.525 177.480 15.805 ;
        RECT 178.985 15.525 179.265 15.805 ;
        RECT 181.840 15.525 182.120 15.805 ;
        RECT 183.625 15.525 183.905 15.805 ;
        RECT 186.480 15.525 186.760 15.805 ;
        RECT 188.265 15.525 188.545 15.805 ;
        RECT 191.120 15.525 191.400 15.805 ;
        RECT 192.905 15.525 193.185 15.805 ;
        RECT 177.200 14.865 177.480 15.145 ;
        RECT 178.985 14.865 179.265 15.145 ;
        RECT 181.840 14.865 182.120 15.145 ;
        RECT 183.625 14.865 183.905 15.145 ;
        RECT 186.480 14.865 186.760 15.145 ;
        RECT 188.265 14.865 188.545 15.145 ;
        RECT 191.120 14.865 191.400 15.145 ;
        RECT 192.905 14.865 193.185 15.145 ;
        RECT 177.200 14.205 177.480 14.485 ;
        RECT 178.985 14.205 179.265 14.485 ;
        RECT 181.840 14.205 182.120 14.485 ;
        RECT 183.625 14.205 183.905 14.485 ;
        RECT 186.480 14.205 186.760 14.485 ;
        RECT 188.265 14.205 188.545 14.485 ;
        RECT 191.120 14.205 191.400 14.485 ;
        RECT 192.905 14.205 193.185 14.485 ;
        RECT 177.200 13.545 177.480 13.825 ;
        RECT 178.985 13.545 179.265 13.825 ;
        RECT 181.840 13.545 182.120 13.825 ;
        RECT 183.625 13.545 183.905 13.825 ;
        RECT 186.480 13.545 186.760 13.825 ;
        RECT 188.265 13.545 188.545 13.825 ;
        RECT 191.120 13.545 191.400 13.825 ;
        RECT 192.905 13.545 193.185 13.825 ;
        RECT 177.200 12.885 177.480 13.165 ;
        RECT 178.985 12.885 179.265 13.165 ;
        RECT 181.840 12.885 182.120 13.165 ;
        RECT 183.625 12.885 183.905 13.165 ;
        RECT 186.480 12.885 186.760 13.165 ;
        RECT 188.265 12.885 188.545 13.165 ;
        RECT 191.120 12.885 191.400 13.165 ;
        RECT 192.905 12.885 193.185 13.165 ;
        RECT 177.200 12.225 177.480 12.505 ;
        RECT 178.985 12.225 179.265 12.505 ;
        RECT 181.840 12.225 182.120 12.505 ;
        RECT 183.625 12.225 183.905 12.505 ;
        RECT 186.480 12.225 186.760 12.505 ;
        RECT 188.265 12.225 188.545 12.505 ;
        RECT 191.120 12.225 191.400 12.505 ;
        RECT 192.905 12.225 193.185 12.505 ;
        RECT 177.200 11.565 177.480 11.845 ;
        RECT 178.985 11.565 179.265 11.845 ;
        RECT 181.840 11.565 182.120 11.845 ;
        RECT 183.625 11.565 183.905 11.845 ;
        RECT 186.480 11.565 186.760 11.845 ;
        RECT 188.265 11.565 188.545 11.845 ;
        RECT 191.120 11.565 191.400 11.845 ;
        RECT 192.905 11.565 193.185 11.845 ;
        RECT 177.200 10.905 177.480 11.185 ;
        RECT 178.985 10.905 179.265 11.185 ;
        RECT 181.840 10.905 182.120 11.185 ;
        RECT 183.625 10.905 183.905 11.185 ;
        RECT 186.480 10.905 186.760 11.185 ;
        RECT 188.265 10.905 188.545 11.185 ;
        RECT 191.120 10.905 191.400 11.185 ;
        RECT 192.905 10.905 193.185 11.185 ;
        RECT 177.200 10.245 177.480 10.525 ;
        RECT 178.985 10.245 179.265 10.525 ;
        RECT 181.840 10.245 182.120 10.525 ;
        RECT 183.625 10.245 183.905 10.525 ;
        RECT 186.480 10.245 186.760 10.525 ;
        RECT 188.265 10.245 188.545 10.525 ;
        RECT 191.120 10.245 191.400 10.525 ;
        RECT 192.905 10.245 193.185 10.525 ;
        RECT 177.200 9.585 177.480 9.865 ;
        RECT 178.985 9.585 179.265 9.865 ;
        RECT 181.840 9.585 182.120 9.865 ;
        RECT 183.625 9.585 183.905 9.865 ;
        RECT 186.480 9.585 186.760 9.865 ;
        RECT 188.265 9.585 188.545 9.865 ;
        RECT 191.120 9.585 191.400 9.865 ;
        RECT 192.905 9.585 193.185 9.865 ;
        RECT 4.660 8.140 4.940 8.420 ;
        RECT 4.660 7.480 4.940 7.760 ;
        RECT 4.660 6.820 4.940 7.100 ;
        RECT 0.900 4.740 1.180 5.020 ;
        RECT 2.040 4.740 2.320 5.020 ;
        RECT 8.080 4.770 8.360 5.050 ;
        RECT 8.740 4.770 9.020 5.050 ;
        RECT 9.400 4.770 9.680 5.050 ;
        RECT 14.610 4.740 14.890 5.020 ;
        RECT 15.270 4.740 15.550 5.020 ;
        RECT 15.930 4.740 16.210 5.020 ;
        RECT 17.970 4.740 18.250 5.020 ;
        RECT 18.630 4.740 18.910 5.020 ;
        RECT 19.290 4.740 19.570 5.020 ;
        RECT 22.850 8.140 23.130 8.420 ;
        RECT 22.850 7.480 23.130 7.760 ;
        RECT 22.850 6.820 23.130 7.100 ;
        RECT 26.270 4.770 26.550 5.050 ;
        RECT 26.930 4.770 27.210 5.050 ;
        RECT 27.590 4.770 27.870 5.050 ;
        RECT 32.800 4.740 33.080 5.020 ;
        RECT 33.460 4.740 33.740 5.020 ;
        RECT 34.120 4.740 34.400 5.020 ;
        RECT 36.160 4.740 36.440 5.020 ;
        RECT 36.820 4.740 37.100 5.020 ;
        RECT 37.480 4.740 37.760 5.020 ;
        RECT 4.220 3.470 4.500 3.750 ;
        RECT 4.630 2.810 4.910 3.090 ;
        RECT 42.160 8.140 42.440 8.420 ;
        RECT 56.990 8.140 57.270 8.420 ;
        RECT 42.160 7.480 42.440 7.760 ;
        RECT 56.990 7.480 57.270 7.760 ;
        RECT 42.160 6.820 42.440 7.100 ;
        RECT 56.990 6.820 57.270 7.100 ;
        RECT 39.540 4.740 39.820 5.020 ;
        RECT 45.580 4.770 45.860 5.050 ;
        RECT 46.240 4.770 46.520 5.050 ;
        RECT 46.900 4.770 47.180 5.050 ;
        RECT 52.110 4.740 52.390 5.020 ;
        RECT 52.770 4.740 53.050 5.020 ;
        RECT 53.430 4.740 53.710 5.020 ;
        RECT 60.410 4.770 60.690 5.050 ;
        RECT 61.070 4.770 61.350 5.050 ;
        RECT 61.730 4.770 62.010 5.050 ;
        RECT 66.940 4.740 67.220 5.020 ;
        RECT 67.600 4.740 67.880 5.020 ;
        RECT 68.260 4.740 68.540 5.020 ;
        RECT 70.300 4.740 70.580 5.020 ;
        RECT 70.960 4.740 71.240 5.020 ;
        RECT 71.620 4.740 71.900 5.020 ;
        RECT 22.410 3.470 22.690 3.750 ;
        RECT 22.820 2.810 23.100 3.090 ;
        RECT 41.720 3.470 42.000 3.750 ;
        RECT 42.130 2.810 42.410 3.090 ;
        RECT 73.680 4.740 73.960 5.020 ;
        RECT 74.680 4.740 74.960 5.020 ;
        RECT 75.340 4.740 75.620 5.020 ;
        RECT 76.000 4.740 76.280 5.020 ;
        RECT 76.920 4.740 77.200 5.020 ;
        RECT 77.580 4.740 77.860 5.020 ;
        RECT 78.240 4.740 78.520 5.020 ;
        RECT 79.260 4.740 79.540 5.020 ;
        RECT 79.920 4.740 80.200 5.020 ;
        RECT 80.580 4.740 80.860 5.020 ;
        RECT 82.520 4.740 82.800 5.020 ;
        RECT 83.180 4.740 83.460 5.020 ;
        RECT 83.840 4.740 84.120 5.020 ;
        RECT 84.760 4.740 85.040 5.020 ;
        RECT 85.420 4.740 85.700 5.020 ;
        RECT 86.080 4.740 86.360 5.020 ;
        RECT 87.000 4.740 87.280 5.020 ;
        RECT 87.660 4.740 87.940 5.020 ;
        RECT 88.320 4.740 88.600 5.020 ;
        RECT 89.240 4.740 89.520 5.020 ;
        RECT 89.900 4.740 90.180 5.020 ;
        RECT 90.560 4.740 90.840 5.020 ;
        RECT 91.480 4.740 91.760 5.020 ;
        RECT 92.140 4.740 92.420 5.020 ;
        RECT 92.800 4.740 93.080 5.020 ;
        RECT 93.840 4.740 94.120 5.020 ;
        RECT 94.840 4.740 95.120 5.020 ;
        RECT 95.500 4.740 95.780 5.020 ;
        RECT 96.160 4.740 96.440 5.020 ;
        RECT 97.080 4.740 97.360 5.020 ;
        RECT 97.740 4.740 98.020 5.020 ;
        RECT 98.400 4.740 98.680 5.020 ;
        RECT 99.320 4.740 99.600 5.020 ;
        RECT 99.980 4.740 100.260 5.020 ;
        RECT 100.640 4.740 100.920 5.020 ;
        RECT 101.660 4.740 101.940 5.020 ;
        RECT 102.320 4.740 102.600 5.020 ;
        RECT 102.980 4.740 103.260 5.020 ;
        RECT 104.920 4.740 105.200 5.020 ;
        RECT 105.580 4.740 105.860 5.020 ;
        RECT 106.240 4.740 106.520 5.020 ;
        RECT 107.160 4.740 107.440 5.020 ;
        RECT 107.820 4.740 108.100 5.020 ;
        RECT 108.480 4.740 108.760 5.020 ;
        RECT 109.400 4.740 109.680 5.020 ;
        RECT 110.060 4.740 110.340 5.020 ;
        RECT 110.720 4.740 111.000 5.020 ;
        RECT 111.640 4.740 111.920 5.020 ;
        RECT 112.300 4.740 112.580 5.020 ;
        RECT 112.960 4.740 113.240 5.020 ;
        RECT 114.000 4.740 114.280 5.020 ;
        RECT 115.000 4.740 115.280 5.020 ;
        RECT 115.660 4.740 115.940 5.020 ;
        RECT 116.320 4.740 116.600 5.020 ;
        RECT 117.240 4.740 117.520 5.020 ;
        RECT 117.900 4.740 118.180 5.020 ;
        RECT 118.560 4.740 118.840 5.020 ;
        RECT 119.480 4.740 119.760 5.020 ;
        RECT 120.140 4.740 120.420 5.020 ;
        RECT 120.800 4.740 121.080 5.020 ;
        RECT 121.820 4.740 122.100 5.020 ;
        RECT 122.480 4.740 122.760 5.020 ;
        RECT 123.140 4.740 123.420 5.020 ;
        RECT 125.080 4.740 125.360 5.020 ;
        RECT 125.740 4.740 126.020 5.020 ;
        RECT 126.400 4.740 126.680 5.020 ;
        RECT 127.320 4.740 127.600 5.020 ;
        RECT 127.980 4.740 128.260 5.020 ;
        RECT 128.640 4.740 128.920 5.020 ;
        RECT 129.560 4.740 129.840 5.020 ;
        RECT 130.220 4.740 130.500 5.020 ;
        RECT 130.880 4.740 131.160 5.020 ;
        RECT 131.800 4.740 132.080 5.020 ;
        RECT 132.460 4.740 132.740 5.020 ;
        RECT 133.120 4.740 133.400 5.020 ;
        RECT 134.160 4.740 134.440 5.020 ;
        RECT 135.160 4.740 135.440 5.020 ;
        RECT 135.820 4.740 136.100 5.020 ;
        RECT 136.480 4.740 136.760 5.020 ;
        RECT 137.400 4.740 137.680 5.020 ;
        RECT 138.060 4.740 138.340 5.020 ;
        RECT 138.720 4.740 139.000 5.020 ;
        RECT 139.640 4.740 139.920 5.020 ;
        RECT 140.300 4.740 140.580 5.020 ;
        RECT 140.960 4.740 141.240 5.020 ;
        RECT 141.880 4.740 142.160 5.020 ;
        RECT 142.540 4.740 142.820 5.020 ;
        RECT 143.200 4.740 143.480 5.020 ;
        RECT 144.220 4.740 144.500 5.020 ;
        RECT 144.880 4.740 145.160 5.020 ;
        RECT 145.540 4.740 145.820 5.020 ;
        RECT 177.200 8.925 177.480 9.205 ;
        RECT 178.985 8.925 179.265 9.205 ;
        RECT 181.840 8.925 182.120 9.205 ;
        RECT 183.625 8.925 183.905 9.205 ;
        RECT 186.480 8.925 186.760 9.205 ;
        RECT 188.265 8.925 188.545 9.205 ;
        RECT 191.120 8.925 191.400 9.205 ;
        RECT 192.905 8.925 193.185 9.205 ;
        RECT 147.480 4.740 147.760 5.020 ;
        RECT 148.140 4.740 148.420 5.020 ;
        RECT 148.800 4.740 149.080 5.020 ;
        RECT 149.720 4.740 150.000 5.020 ;
        RECT 150.380 4.740 150.660 5.020 ;
        RECT 151.040 4.740 151.320 5.020 ;
        RECT 151.960 4.740 152.240 5.020 ;
        RECT 152.620 4.740 152.900 5.020 ;
        RECT 153.280 4.740 153.560 5.020 ;
        RECT 154.320 4.740 154.600 5.020 ;
        RECT 155.320 4.740 155.600 5.020 ;
        RECT 155.980 4.740 156.260 5.020 ;
        RECT 156.640 4.740 156.920 5.020 ;
        RECT 157.560 4.740 157.840 5.020 ;
        RECT 158.220 4.740 158.500 5.020 ;
        RECT 158.880 4.740 159.160 5.020 ;
        RECT 159.800 4.740 160.080 5.020 ;
        RECT 160.460 4.740 160.740 5.020 ;
        RECT 161.120 4.740 161.400 5.020 ;
        RECT 162.040 4.740 162.320 5.020 ;
        RECT 162.700 4.740 162.980 5.020 ;
        RECT 163.360 4.740 163.640 5.020 ;
        RECT 164.280 4.740 164.560 5.020 ;
        RECT 164.940 4.740 165.220 5.020 ;
        RECT 165.600 4.740 165.880 5.020 ;
        RECT 166.620 4.740 166.900 5.020 ;
        RECT 167.280 4.740 167.560 5.020 ;
        RECT 167.940 4.740 168.220 5.020 ;
        RECT 169.880 4.740 170.160 5.020 ;
        RECT 170.540 4.740 170.820 5.020 ;
        RECT 171.200 4.740 171.480 5.020 ;
        RECT 172.120 4.740 172.400 5.020 ;
        RECT 172.780 4.740 173.060 5.020 ;
        RECT 173.440 4.740 173.720 5.020 ;
        RECT 174.460 4.740 174.740 5.020 ;
        RECT 56.550 3.470 56.830 3.750 ;
        RECT 56.960 2.810 57.240 3.090 ;
        RECT 0.900 0.820 1.180 1.100 ;
        RECT 2.040 0.820 2.320 1.100 ;
        RECT 7.480 0.820 7.760 1.100 ;
        RECT 8.140 0.820 8.420 1.100 ;
        RECT 8.800 0.820 9.080 1.100 ;
        RECT 14.350 0.820 14.630 1.100 ;
        RECT 15.670 0.820 15.950 1.100 ;
        RECT 17.710 0.820 17.990 1.100 ;
        RECT 19.030 0.820 19.310 1.100 ;
        RECT 25.670 0.820 25.950 1.100 ;
        RECT 26.330 0.820 26.610 1.100 ;
        RECT 26.990 0.820 27.270 1.100 ;
        RECT 32.540 0.820 32.820 1.100 ;
        RECT 33.860 0.820 34.140 1.100 ;
        RECT 35.900 0.820 36.180 1.100 ;
        RECT 37.220 0.820 37.500 1.100 ;
        RECT 39.540 0.820 39.820 1.100 ;
        RECT 44.980 0.820 45.260 1.100 ;
        RECT 45.640 0.820 45.920 1.100 ;
        RECT 46.300 0.820 46.580 1.100 ;
        RECT 51.850 0.820 52.130 1.100 ;
        RECT 53.170 0.820 53.450 1.100 ;
        RECT 59.810 0.820 60.090 1.100 ;
        RECT 60.470 0.820 60.750 1.100 ;
        RECT 61.130 0.820 61.410 1.100 ;
        RECT 66.680 0.820 66.960 1.100 ;
        RECT 68.000 0.820 68.280 1.100 ;
        RECT 70.040 0.820 70.320 1.100 ;
        RECT 71.360 0.820 71.640 1.100 ;
        RECT 73.680 0.820 73.960 1.100 ;
        RECT 74.680 0.820 74.960 1.100 ;
        RECT 75.340 0.820 75.620 1.100 ;
        RECT 76.000 0.820 76.280 1.100 ;
        RECT 76.920 0.820 77.200 1.100 ;
        RECT 77.580 0.820 77.860 1.100 ;
        RECT 78.240 0.820 78.520 1.100 ;
        RECT 79.000 0.820 79.280 1.100 ;
        RECT 80.320 0.820 80.600 1.100 ;
        RECT 82.520 0.820 82.800 1.100 ;
        RECT 83.180 0.820 83.460 1.100 ;
        RECT 83.840 0.820 84.120 1.100 ;
        RECT 84.760 0.820 85.040 1.100 ;
        RECT 85.420 0.820 85.700 1.100 ;
        RECT 86.080 0.820 86.360 1.100 ;
        RECT 87.000 0.820 87.280 1.100 ;
        RECT 87.660 0.820 87.940 1.100 ;
        RECT 88.320 0.820 88.600 1.100 ;
        RECT 89.240 0.820 89.520 1.100 ;
        RECT 89.900 0.820 90.180 1.100 ;
        RECT 90.560 0.820 90.840 1.100 ;
        RECT 91.480 0.820 91.760 1.100 ;
        RECT 92.140 0.820 92.420 1.100 ;
        RECT 92.800 0.820 93.080 1.100 ;
        RECT 93.840 0.820 94.120 1.100 ;
        RECT 94.840 0.820 95.120 1.100 ;
        RECT 95.500 0.820 95.780 1.100 ;
        RECT 96.160 0.820 96.440 1.100 ;
        RECT 97.080 0.820 97.360 1.100 ;
        RECT 97.740 0.820 98.020 1.100 ;
        RECT 98.400 0.820 98.680 1.100 ;
        RECT 99.320 0.820 99.600 1.100 ;
        RECT 99.980 0.820 100.260 1.100 ;
        RECT 100.640 0.820 100.920 1.100 ;
        RECT 101.400 0.820 101.680 1.100 ;
        RECT 102.720 0.820 103.000 1.100 ;
        RECT 104.920 0.820 105.200 1.100 ;
        RECT 105.580 0.820 105.860 1.100 ;
        RECT 106.240 0.820 106.520 1.100 ;
        RECT 107.160 0.820 107.440 1.100 ;
        RECT 107.820 0.820 108.100 1.100 ;
        RECT 108.480 0.820 108.760 1.100 ;
        RECT 109.400 0.820 109.680 1.100 ;
        RECT 110.060 0.820 110.340 1.100 ;
        RECT 110.720 0.820 111.000 1.100 ;
        RECT 111.640 0.820 111.920 1.100 ;
        RECT 112.300 0.820 112.580 1.100 ;
        RECT 112.960 0.820 113.240 1.100 ;
        RECT 114.000 0.820 114.280 1.100 ;
        RECT 115.000 0.820 115.280 1.100 ;
        RECT 115.660 0.820 115.940 1.100 ;
        RECT 116.320 0.820 116.600 1.100 ;
        RECT 117.240 0.820 117.520 1.100 ;
        RECT 117.900 0.820 118.180 1.100 ;
        RECT 118.560 0.820 118.840 1.100 ;
        RECT 119.480 0.820 119.760 1.100 ;
        RECT 120.140 0.820 120.420 1.100 ;
        RECT 120.800 0.820 121.080 1.100 ;
        RECT 121.560 0.820 121.840 1.100 ;
        RECT 122.880 0.820 123.160 1.100 ;
        RECT 125.080 0.820 125.360 1.100 ;
        RECT 125.740 0.820 126.020 1.100 ;
        RECT 126.400 0.820 126.680 1.100 ;
        RECT 127.320 0.820 127.600 1.100 ;
        RECT 127.980 0.820 128.260 1.100 ;
        RECT 128.640 0.820 128.920 1.100 ;
        RECT 129.560 0.820 129.840 1.100 ;
        RECT 130.220 0.820 130.500 1.100 ;
        RECT 130.880 0.820 131.160 1.100 ;
        RECT 131.800 0.820 132.080 1.100 ;
        RECT 132.460 0.820 132.740 1.100 ;
        RECT 133.120 0.820 133.400 1.100 ;
        RECT 134.160 0.820 134.440 1.100 ;
        RECT 135.160 0.820 135.440 1.100 ;
        RECT 135.820 0.820 136.100 1.100 ;
        RECT 136.480 0.820 136.760 1.100 ;
        RECT 137.400 0.820 137.680 1.100 ;
        RECT 138.060 0.820 138.340 1.100 ;
        RECT 138.720 0.820 139.000 1.100 ;
        RECT 139.640 0.820 139.920 1.100 ;
        RECT 140.300 0.820 140.580 1.100 ;
        RECT 140.960 0.820 141.240 1.100 ;
        RECT 141.880 0.820 142.160 1.100 ;
        RECT 142.540 0.820 142.820 1.100 ;
        RECT 143.200 0.820 143.480 1.100 ;
        RECT 143.960 0.820 144.240 1.100 ;
        RECT 145.280 0.820 145.560 1.100 ;
        RECT 147.480 0.820 147.760 1.100 ;
        RECT 148.140 0.820 148.420 1.100 ;
        RECT 148.800 0.820 149.080 1.100 ;
        RECT 149.720 0.820 150.000 1.100 ;
        RECT 150.380 0.820 150.660 1.100 ;
        RECT 151.040 0.820 151.320 1.100 ;
        RECT 151.960 0.820 152.240 1.100 ;
        RECT 152.620 0.820 152.900 1.100 ;
        RECT 153.280 0.820 153.560 1.100 ;
        RECT 154.320 0.820 154.600 1.100 ;
        RECT 155.320 0.820 155.600 1.100 ;
        RECT 155.980 0.820 156.260 1.100 ;
        RECT 156.640 0.820 156.920 1.100 ;
        RECT 157.560 0.820 157.840 1.100 ;
        RECT 158.220 0.820 158.500 1.100 ;
        RECT 158.880 0.820 159.160 1.100 ;
        RECT 159.800 0.820 160.080 1.100 ;
        RECT 160.460 0.820 160.740 1.100 ;
        RECT 161.120 0.820 161.400 1.100 ;
        RECT 162.040 0.820 162.320 1.100 ;
        RECT 162.700 0.820 162.980 1.100 ;
        RECT 163.360 0.820 163.640 1.100 ;
        RECT 164.280 0.820 164.560 1.100 ;
        RECT 164.940 0.820 165.220 1.100 ;
        RECT 165.600 0.820 165.880 1.100 ;
        RECT 166.360 0.820 166.640 1.100 ;
        RECT 167.680 0.820 167.960 1.100 ;
        RECT 169.880 0.820 170.160 1.100 ;
        RECT 170.540 0.820 170.820 1.100 ;
        RECT 171.200 0.820 171.480 1.100 ;
        RECT 172.120 0.820 172.400 1.100 ;
        RECT 172.780 0.820 173.060 1.100 ;
        RECT 173.440 0.820 173.720 1.100 ;
        RECT 174.460 0.820 174.740 1.100 ;
      LAYER Metal3 ;
        RECT 0.765 58.745 1.145 59.125 ;
        RECT 11.055 58.745 11.435 59.125 ;
        RECT 21.340 58.745 21.720 59.125 ;
        RECT 22.760 58.745 23.140 59.125 ;
        RECT 33.050 58.745 33.430 59.125 ;
        RECT 43.335 58.745 43.715 59.125 ;
        RECT 44.755 58.745 45.135 59.125 ;
        RECT 55.045 58.745 55.425 59.125 ;
        RECT 65.330 58.745 65.710 59.125 ;
        RECT 66.750 58.745 67.130 59.125 ;
        RECT 77.040 58.745 77.420 59.125 ;
        RECT 87.325 58.745 87.705 59.125 ;
        RECT 88.745 58.745 89.125 59.125 ;
        RECT 99.035 58.745 99.415 59.125 ;
        RECT 109.320 58.745 109.700 59.125 ;
        RECT 110.740 58.745 111.120 59.125 ;
        RECT 121.030 58.745 121.410 59.125 ;
        RECT 131.315 58.745 131.695 59.125 ;
        RECT 132.735 58.745 133.115 59.125 ;
        RECT 143.025 58.745 143.405 59.125 ;
        RECT 153.310 58.745 153.690 59.125 ;
        RECT 154.730 58.745 155.110 59.125 ;
        RECT 165.020 58.745 165.400 59.125 ;
        RECT 175.305 58.745 175.685 59.125 ;
        RECT 0.765 58.085 1.145 58.465 ;
        RECT 11.055 58.085 11.435 58.465 ;
        RECT 21.340 58.085 21.720 58.465 ;
        RECT 22.760 58.085 23.140 58.465 ;
        RECT 33.050 58.085 33.430 58.465 ;
        RECT 43.335 58.085 43.715 58.465 ;
        RECT 44.755 58.085 45.135 58.465 ;
        RECT 55.045 58.085 55.425 58.465 ;
        RECT 65.330 58.085 65.710 58.465 ;
        RECT 66.750 58.085 67.130 58.465 ;
        RECT 77.040 58.085 77.420 58.465 ;
        RECT 87.325 58.085 87.705 58.465 ;
        RECT 88.745 58.085 89.125 58.465 ;
        RECT 99.035 58.085 99.415 58.465 ;
        RECT 109.320 58.085 109.700 58.465 ;
        RECT 110.740 58.085 111.120 58.465 ;
        RECT 121.030 58.085 121.410 58.465 ;
        RECT 131.315 58.085 131.695 58.465 ;
        RECT 132.735 58.085 133.115 58.465 ;
        RECT 143.025 58.085 143.405 58.465 ;
        RECT 153.310 58.085 153.690 58.465 ;
        RECT 154.730 58.085 155.110 58.465 ;
        RECT 165.020 58.085 165.400 58.465 ;
        RECT 175.305 58.085 175.685 58.465 ;
        RECT 0.765 57.425 1.145 57.805 ;
        RECT 11.055 57.425 11.435 57.805 ;
        RECT 21.340 57.425 21.720 57.805 ;
        RECT 22.760 57.425 23.140 57.805 ;
        RECT 33.050 57.425 33.430 57.805 ;
        RECT 43.335 57.425 43.715 57.805 ;
        RECT 44.755 57.425 45.135 57.805 ;
        RECT 55.045 57.425 55.425 57.805 ;
        RECT 65.330 57.425 65.710 57.805 ;
        RECT 66.750 57.425 67.130 57.805 ;
        RECT 77.040 57.425 77.420 57.805 ;
        RECT 87.325 57.425 87.705 57.805 ;
        RECT 88.745 57.425 89.125 57.805 ;
        RECT 99.035 57.425 99.415 57.805 ;
        RECT 109.320 57.425 109.700 57.805 ;
        RECT 110.740 57.425 111.120 57.805 ;
        RECT 121.030 57.425 121.410 57.805 ;
        RECT 131.315 57.425 131.695 57.805 ;
        RECT 132.735 57.425 133.115 57.805 ;
        RECT 143.025 57.425 143.405 57.805 ;
        RECT 153.310 57.425 153.690 57.805 ;
        RECT 154.730 57.425 155.110 57.805 ;
        RECT 165.020 57.425 165.400 57.805 ;
        RECT 175.305 57.425 175.685 57.805 ;
        RECT 0.765 56.765 1.145 57.145 ;
        RECT 11.055 56.765 11.435 57.145 ;
        RECT 21.340 56.765 21.720 57.145 ;
        RECT 22.760 56.765 23.140 57.145 ;
        RECT 33.050 56.765 33.430 57.145 ;
        RECT 43.335 56.765 43.715 57.145 ;
        RECT 44.755 56.765 45.135 57.145 ;
        RECT 55.045 56.765 55.425 57.145 ;
        RECT 65.330 56.765 65.710 57.145 ;
        RECT 66.750 56.765 67.130 57.145 ;
        RECT 77.040 56.765 77.420 57.145 ;
        RECT 87.325 56.765 87.705 57.145 ;
        RECT 88.745 56.765 89.125 57.145 ;
        RECT 99.035 56.765 99.415 57.145 ;
        RECT 109.320 56.765 109.700 57.145 ;
        RECT 110.740 56.765 111.120 57.145 ;
        RECT 121.030 56.765 121.410 57.145 ;
        RECT 131.315 56.765 131.695 57.145 ;
        RECT 132.735 56.765 133.115 57.145 ;
        RECT 143.025 56.765 143.405 57.145 ;
        RECT 153.310 56.765 153.690 57.145 ;
        RECT 154.730 56.765 155.110 57.145 ;
        RECT 165.020 56.765 165.400 57.145 ;
        RECT 175.305 56.765 175.685 57.145 ;
        RECT 0.765 56.105 1.145 56.485 ;
        RECT 11.055 56.105 11.435 56.485 ;
        RECT 21.340 56.105 21.720 56.485 ;
        RECT 22.760 56.105 23.140 56.485 ;
        RECT 33.050 56.105 33.430 56.485 ;
        RECT 43.335 56.105 43.715 56.485 ;
        RECT 44.755 56.105 45.135 56.485 ;
        RECT 55.045 56.105 55.425 56.485 ;
        RECT 65.330 56.105 65.710 56.485 ;
        RECT 66.750 56.105 67.130 56.485 ;
        RECT 77.040 56.105 77.420 56.485 ;
        RECT 87.325 56.105 87.705 56.485 ;
        RECT 88.745 56.105 89.125 56.485 ;
        RECT 99.035 56.105 99.415 56.485 ;
        RECT 109.320 56.105 109.700 56.485 ;
        RECT 110.740 56.105 111.120 56.485 ;
        RECT 121.030 56.105 121.410 56.485 ;
        RECT 131.315 56.105 131.695 56.485 ;
        RECT 132.735 56.105 133.115 56.485 ;
        RECT 143.025 56.105 143.405 56.485 ;
        RECT 153.310 56.105 153.690 56.485 ;
        RECT 154.730 56.105 155.110 56.485 ;
        RECT 165.020 56.105 165.400 56.485 ;
        RECT 175.305 56.105 175.685 56.485 ;
        RECT 0.765 55.445 1.145 55.825 ;
        RECT 11.055 55.445 11.435 55.825 ;
        RECT 21.340 55.445 21.720 55.825 ;
        RECT 22.760 55.445 23.140 55.825 ;
        RECT 33.050 55.445 33.430 55.825 ;
        RECT 43.335 55.445 43.715 55.825 ;
        RECT 44.755 55.445 45.135 55.825 ;
        RECT 55.045 55.445 55.425 55.825 ;
        RECT 65.330 55.445 65.710 55.825 ;
        RECT 66.750 55.445 67.130 55.825 ;
        RECT 77.040 55.445 77.420 55.825 ;
        RECT 87.325 55.445 87.705 55.825 ;
        RECT 88.745 55.445 89.125 55.825 ;
        RECT 99.035 55.445 99.415 55.825 ;
        RECT 109.320 55.445 109.700 55.825 ;
        RECT 110.740 55.445 111.120 55.825 ;
        RECT 121.030 55.445 121.410 55.825 ;
        RECT 131.315 55.445 131.695 55.825 ;
        RECT 132.735 55.445 133.115 55.825 ;
        RECT 143.025 55.445 143.405 55.825 ;
        RECT 153.310 55.445 153.690 55.825 ;
        RECT 154.730 55.445 155.110 55.825 ;
        RECT 165.020 55.445 165.400 55.825 ;
        RECT 175.305 55.445 175.685 55.825 ;
        RECT 0.765 54.785 1.145 55.165 ;
        RECT 11.055 54.785 11.435 55.165 ;
        RECT 21.340 54.785 21.720 55.165 ;
        RECT 22.760 54.785 23.140 55.165 ;
        RECT 33.050 54.785 33.430 55.165 ;
        RECT 43.335 54.785 43.715 55.165 ;
        RECT 44.755 54.785 45.135 55.165 ;
        RECT 55.045 54.785 55.425 55.165 ;
        RECT 65.330 54.785 65.710 55.165 ;
        RECT 66.750 54.785 67.130 55.165 ;
        RECT 77.040 54.785 77.420 55.165 ;
        RECT 87.325 54.785 87.705 55.165 ;
        RECT 88.745 54.785 89.125 55.165 ;
        RECT 99.035 54.785 99.415 55.165 ;
        RECT 109.320 54.785 109.700 55.165 ;
        RECT 110.740 54.785 111.120 55.165 ;
        RECT 121.030 54.785 121.410 55.165 ;
        RECT 131.315 54.785 131.695 55.165 ;
        RECT 132.735 54.785 133.115 55.165 ;
        RECT 143.025 54.785 143.405 55.165 ;
        RECT 153.310 54.785 153.690 55.165 ;
        RECT 154.730 54.785 155.110 55.165 ;
        RECT 165.020 54.785 165.400 55.165 ;
        RECT 175.305 54.785 175.685 55.165 ;
        RECT 177.150 55.115 177.530 55.495 ;
        RECT 178.935 55.115 179.315 55.495 ;
        RECT 181.790 55.115 182.170 55.495 ;
        RECT 183.575 55.115 183.955 55.495 ;
        RECT 186.430 55.115 186.810 55.495 ;
        RECT 188.215 55.115 188.595 55.495 ;
        RECT 191.070 55.115 191.450 55.495 ;
        RECT 192.855 55.115 193.235 55.495 ;
        RECT 0.765 54.125 1.145 54.505 ;
        RECT 11.055 54.125 11.435 54.505 ;
        RECT 21.340 54.125 21.720 54.505 ;
        RECT 22.760 54.125 23.140 54.505 ;
        RECT 33.050 54.125 33.430 54.505 ;
        RECT 43.335 54.125 43.715 54.505 ;
        RECT 44.755 54.125 45.135 54.505 ;
        RECT 55.045 54.125 55.425 54.505 ;
        RECT 65.330 54.125 65.710 54.505 ;
        RECT 66.750 54.125 67.130 54.505 ;
        RECT 77.040 54.125 77.420 54.505 ;
        RECT 87.325 54.125 87.705 54.505 ;
        RECT 88.745 54.125 89.125 54.505 ;
        RECT 99.035 54.125 99.415 54.505 ;
        RECT 109.320 54.125 109.700 54.505 ;
        RECT 110.740 54.125 111.120 54.505 ;
        RECT 121.030 54.125 121.410 54.505 ;
        RECT 131.315 54.125 131.695 54.505 ;
        RECT 132.735 54.125 133.115 54.505 ;
        RECT 143.025 54.125 143.405 54.505 ;
        RECT 153.310 54.125 153.690 54.505 ;
        RECT 154.730 54.125 155.110 54.505 ;
        RECT 165.020 54.125 165.400 54.505 ;
        RECT 175.305 54.125 175.685 54.505 ;
        RECT 177.150 54.455 177.530 54.835 ;
        RECT 178.935 54.455 179.315 54.835 ;
        RECT 181.790 54.455 182.170 54.835 ;
        RECT 183.575 54.455 183.955 54.835 ;
        RECT 186.430 54.455 186.810 54.835 ;
        RECT 188.215 54.455 188.595 54.835 ;
        RECT 191.070 54.455 191.450 54.835 ;
        RECT 192.855 54.455 193.235 54.835 ;
        RECT 0.765 53.465 1.145 53.845 ;
        RECT 11.055 53.465 11.435 53.845 ;
        RECT 21.340 53.465 21.720 53.845 ;
        RECT 22.760 53.465 23.140 53.845 ;
        RECT 33.050 53.465 33.430 53.845 ;
        RECT 43.335 53.465 43.715 53.845 ;
        RECT 44.755 53.465 45.135 53.845 ;
        RECT 55.045 53.465 55.425 53.845 ;
        RECT 65.330 53.465 65.710 53.845 ;
        RECT 66.750 53.465 67.130 53.845 ;
        RECT 77.040 53.465 77.420 53.845 ;
        RECT 87.325 53.465 87.705 53.845 ;
        RECT 88.745 53.465 89.125 53.845 ;
        RECT 99.035 53.465 99.415 53.845 ;
        RECT 109.320 53.465 109.700 53.845 ;
        RECT 110.740 53.465 111.120 53.845 ;
        RECT 121.030 53.465 121.410 53.845 ;
        RECT 131.315 53.465 131.695 53.845 ;
        RECT 132.735 53.465 133.115 53.845 ;
        RECT 143.025 53.465 143.405 53.845 ;
        RECT 153.310 53.465 153.690 53.845 ;
        RECT 154.730 53.465 155.110 53.845 ;
        RECT 165.020 53.465 165.400 53.845 ;
        RECT 175.305 53.465 175.685 53.845 ;
        RECT 177.150 53.795 177.530 54.175 ;
        RECT 178.935 53.795 179.315 54.175 ;
        RECT 181.790 53.795 182.170 54.175 ;
        RECT 183.575 53.795 183.955 54.175 ;
        RECT 186.430 53.795 186.810 54.175 ;
        RECT 188.215 53.795 188.595 54.175 ;
        RECT 191.070 53.795 191.450 54.175 ;
        RECT 192.855 53.795 193.235 54.175 ;
        RECT 0.765 52.805 1.145 53.185 ;
        RECT 11.055 52.805 11.435 53.185 ;
        RECT 21.340 52.805 21.720 53.185 ;
        RECT 22.760 52.805 23.140 53.185 ;
        RECT 33.050 52.805 33.430 53.185 ;
        RECT 43.335 52.805 43.715 53.185 ;
        RECT 44.755 52.805 45.135 53.185 ;
        RECT 55.045 52.805 55.425 53.185 ;
        RECT 65.330 52.805 65.710 53.185 ;
        RECT 66.750 52.805 67.130 53.185 ;
        RECT 77.040 52.805 77.420 53.185 ;
        RECT 87.325 52.805 87.705 53.185 ;
        RECT 88.745 52.805 89.125 53.185 ;
        RECT 99.035 52.805 99.415 53.185 ;
        RECT 109.320 52.805 109.700 53.185 ;
        RECT 110.740 52.805 111.120 53.185 ;
        RECT 121.030 52.805 121.410 53.185 ;
        RECT 131.315 52.805 131.695 53.185 ;
        RECT 132.735 52.805 133.115 53.185 ;
        RECT 143.025 52.805 143.405 53.185 ;
        RECT 153.310 52.805 153.690 53.185 ;
        RECT 154.730 52.805 155.110 53.185 ;
        RECT 165.020 52.805 165.400 53.185 ;
        RECT 175.305 52.805 175.685 53.185 ;
        RECT 177.150 53.135 177.530 53.515 ;
        RECT 178.935 53.135 179.315 53.515 ;
        RECT 181.790 53.135 182.170 53.515 ;
        RECT 183.575 53.135 183.955 53.515 ;
        RECT 186.430 53.135 186.810 53.515 ;
        RECT 188.215 53.135 188.595 53.515 ;
        RECT 191.070 53.135 191.450 53.515 ;
        RECT 192.855 53.135 193.235 53.515 ;
        RECT 0.765 52.145 1.145 52.525 ;
        RECT 11.055 52.145 11.435 52.525 ;
        RECT 21.340 52.145 21.720 52.525 ;
        RECT 22.760 52.145 23.140 52.525 ;
        RECT 33.050 52.145 33.430 52.525 ;
        RECT 43.335 52.145 43.715 52.525 ;
        RECT 44.755 52.145 45.135 52.525 ;
        RECT 55.045 52.145 55.425 52.525 ;
        RECT 65.330 52.145 65.710 52.525 ;
        RECT 66.750 52.145 67.130 52.525 ;
        RECT 77.040 52.145 77.420 52.525 ;
        RECT 87.325 52.145 87.705 52.525 ;
        RECT 88.745 52.145 89.125 52.525 ;
        RECT 99.035 52.145 99.415 52.525 ;
        RECT 109.320 52.145 109.700 52.525 ;
        RECT 110.740 52.145 111.120 52.525 ;
        RECT 121.030 52.145 121.410 52.525 ;
        RECT 131.315 52.145 131.695 52.525 ;
        RECT 132.735 52.145 133.115 52.525 ;
        RECT 143.025 52.145 143.405 52.525 ;
        RECT 153.310 52.145 153.690 52.525 ;
        RECT 154.730 52.145 155.110 52.525 ;
        RECT 165.020 52.145 165.400 52.525 ;
        RECT 175.305 52.145 175.685 52.525 ;
        RECT 177.150 52.475 177.530 52.855 ;
        RECT 178.935 52.475 179.315 52.855 ;
        RECT 181.790 52.475 182.170 52.855 ;
        RECT 183.575 52.475 183.955 52.855 ;
        RECT 186.430 52.475 186.810 52.855 ;
        RECT 188.215 52.475 188.595 52.855 ;
        RECT 191.070 52.475 191.450 52.855 ;
        RECT 192.855 52.475 193.235 52.855 ;
        RECT 0.765 51.485 1.145 51.865 ;
        RECT 11.055 51.485 11.435 51.865 ;
        RECT 21.340 51.485 21.720 51.865 ;
        RECT 22.760 51.485 23.140 51.865 ;
        RECT 33.050 51.485 33.430 51.865 ;
        RECT 43.335 51.485 43.715 51.865 ;
        RECT 44.755 51.485 45.135 51.865 ;
        RECT 55.045 51.485 55.425 51.865 ;
        RECT 65.330 51.485 65.710 51.865 ;
        RECT 66.750 51.485 67.130 51.865 ;
        RECT 77.040 51.485 77.420 51.865 ;
        RECT 87.325 51.485 87.705 51.865 ;
        RECT 88.745 51.485 89.125 51.865 ;
        RECT 99.035 51.485 99.415 51.865 ;
        RECT 109.320 51.485 109.700 51.865 ;
        RECT 110.740 51.485 111.120 51.865 ;
        RECT 121.030 51.485 121.410 51.865 ;
        RECT 131.315 51.485 131.695 51.865 ;
        RECT 132.735 51.485 133.115 51.865 ;
        RECT 143.025 51.485 143.405 51.865 ;
        RECT 153.310 51.485 153.690 51.865 ;
        RECT 154.730 51.485 155.110 51.865 ;
        RECT 165.020 51.485 165.400 51.865 ;
        RECT 175.305 51.485 175.685 51.865 ;
        RECT 177.150 51.815 177.530 52.195 ;
        RECT 178.935 51.815 179.315 52.195 ;
        RECT 181.790 51.815 182.170 52.195 ;
        RECT 183.575 51.815 183.955 52.195 ;
        RECT 186.430 51.815 186.810 52.195 ;
        RECT 188.215 51.815 188.595 52.195 ;
        RECT 191.070 51.815 191.450 52.195 ;
        RECT 192.855 51.815 193.235 52.195 ;
        RECT 0.765 50.825 1.145 51.205 ;
        RECT 11.055 50.825 11.435 51.205 ;
        RECT 21.340 50.825 21.720 51.205 ;
        RECT 22.760 50.825 23.140 51.205 ;
        RECT 33.050 50.825 33.430 51.205 ;
        RECT 43.335 50.825 43.715 51.205 ;
        RECT 44.755 50.825 45.135 51.205 ;
        RECT 55.045 50.825 55.425 51.205 ;
        RECT 65.330 50.825 65.710 51.205 ;
        RECT 66.750 50.825 67.130 51.205 ;
        RECT 77.040 50.825 77.420 51.205 ;
        RECT 87.325 50.825 87.705 51.205 ;
        RECT 88.745 50.825 89.125 51.205 ;
        RECT 99.035 50.825 99.415 51.205 ;
        RECT 109.320 50.825 109.700 51.205 ;
        RECT 110.740 50.825 111.120 51.205 ;
        RECT 121.030 50.825 121.410 51.205 ;
        RECT 131.315 50.825 131.695 51.205 ;
        RECT 132.735 50.825 133.115 51.205 ;
        RECT 143.025 50.825 143.405 51.205 ;
        RECT 153.310 50.825 153.690 51.205 ;
        RECT 154.730 50.825 155.110 51.205 ;
        RECT 165.020 50.825 165.400 51.205 ;
        RECT 175.305 50.825 175.685 51.205 ;
        RECT 177.150 51.155 177.530 51.535 ;
        RECT 178.935 51.155 179.315 51.535 ;
        RECT 181.790 51.155 182.170 51.535 ;
        RECT 183.575 51.155 183.955 51.535 ;
        RECT 186.430 51.155 186.810 51.535 ;
        RECT 188.215 51.155 188.595 51.535 ;
        RECT 191.070 51.155 191.450 51.535 ;
        RECT 192.855 51.155 193.235 51.535 ;
        RECT 0.765 50.165 1.145 50.545 ;
        RECT 11.055 50.165 11.435 50.545 ;
        RECT 21.340 50.165 21.720 50.545 ;
        RECT 22.760 50.165 23.140 50.545 ;
        RECT 33.050 50.165 33.430 50.545 ;
        RECT 43.335 50.165 43.715 50.545 ;
        RECT 44.755 50.165 45.135 50.545 ;
        RECT 55.045 50.165 55.425 50.545 ;
        RECT 65.330 50.165 65.710 50.545 ;
        RECT 66.750 50.165 67.130 50.545 ;
        RECT 77.040 50.165 77.420 50.545 ;
        RECT 87.325 50.165 87.705 50.545 ;
        RECT 88.745 50.165 89.125 50.545 ;
        RECT 99.035 50.165 99.415 50.545 ;
        RECT 109.320 50.165 109.700 50.545 ;
        RECT 110.740 50.165 111.120 50.545 ;
        RECT 121.030 50.165 121.410 50.545 ;
        RECT 131.315 50.165 131.695 50.545 ;
        RECT 132.735 50.165 133.115 50.545 ;
        RECT 143.025 50.165 143.405 50.545 ;
        RECT 153.310 50.165 153.690 50.545 ;
        RECT 154.730 50.165 155.110 50.545 ;
        RECT 165.020 50.165 165.400 50.545 ;
        RECT 175.305 50.165 175.685 50.545 ;
        RECT 177.150 50.495 177.530 50.875 ;
        RECT 178.935 50.495 179.315 50.875 ;
        RECT 181.790 50.495 182.170 50.875 ;
        RECT 183.575 50.495 183.955 50.875 ;
        RECT 186.430 50.495 186.810 50.875 ;
        RECT 188.215 50.495 188.595 50.875 ;
        RECT 191.070 50.495 191.450 50.875 ;
        RECT 192.855 50.495 193.235 50.875 ;
        RECT 0.500 46.485 193.820 48.185 ;
        RECT 0.500 43.785 193.820 45.485 ;
        RECT 0.500 23.585 193.820 25.285 ;
        RECT 0.500 20.885 193.820 22.585 ;
        RECT 177.150 18.115 177.530 18.495 ;
        RECT 178.935 18.115 179.315 18.495 ;
        RECT 181.790 18.115 182.170 18.495 ;
        RECT 183.575 18.115 183.955 18.495 ;
        RECT 186.430 18.115 186.810 18.495 ;
        RECT 188.215 18.115 188.595 18.495 ;
        RECT 191.070 18.115 191.450 18.495 ;
        RECT 192.855 18.115 193.235 18.495 ;
        RECT 177.150 17.455 177.530 17.835 ;
        RECT 178.935 17.455 179.315 17.835 ;
        RECT 181.790 17.455 182.170 17.835 ;
        RECT 183.575 17.455 183.955 17.835 ;
        RECT 186.430 17.455 186.810 17.835 ;
        RECT 188.215 17.455 188.595 17.835 ;
        RECT 191.070 17.455 191.450 17.835 ;
        RECT 192.855 17.455 193.235 17.835 ;
        RECT 177.150 16.795 177.530 17.175 ;
        RECT 178.935 16.795 179.315 17.175 ;
        RECT 181.790 16.795 182.170 17.175 ;
        RECT 183.575 16.795 183.955 17.175 ;
        RECT 186.430 16.795 186.810 17.175 ;
        RECT 188.215 16.795 188.595 17.175 ;
        RECT 191.070 16.795 191.450 17.175 ;
        RECT 192.855 16.795 193.235 17.175 ;
        RECT 177.150 16.135 177.530 16.515 ;
        RECT 178.935 16.135 179.315 16.515 ;
        RECT 181.790 16.135 182.170 16.515 ;
        RECT 183.575 16.135 183.955 16.515 ;
        RECT 186.430 16.135 186.810 16.515 ;
        RECT 188.215 16.135 188.595 16.515 ;
        RECT 191.070 16.135 191.450 16.515 ;
        RECT 192.855 16.135 193.235 16.515 ;
        RECT 177.150 15.475 177.530 15.855 ;
        RECT 178.935 15.475 179.315 15.855 ;
        RECT 181.790 15.475 182.170 15.855 ;
        RECT 183.575 15.475 183.955 15.855 ;
        RECT 186.430 15.475 186.810 15.855 ;
        RECT 188.215 15.475 188.595 15.855 ;
        RECT 191.070 15.475 191.450 15.855 ;
        RECT 192.855 15.475 193.235 15.855 ;
        RECT 177.150 14.815 177.530 15.195 ;
        RECT 178.935 14.815 179.315 15.195 ;
        RECT 181.790 14.815 182.170 15.195 ;
        RECT 183.575 14.815 183.955 15.195 ;
        RECT 186.430 14.815 186.810 15.195 ;
        RECT 188.215 14.815 188.595 15.195 ;
        RECT 191.070 14.815 191.450 15.195 ;
        RECT 192.855 14.815 193.235 15.195 ;
        RECT 177.150 14.155 177.530 14.535 ;
        RECT 178.935 14.155 179.315 14.535 ;
        RECT 181.790 14.155 182.170 14.535 ;
        RECT 183.575 14.155 183.955 14.535 ;
        RECT 186.430 14.155 186.810 14.535 ;
        RECT 188.215 14.155 188.595 14.535 ;
        RECT 191.070 14.155 191.450 14.535 ;
        RECT 192.855 14.155 193.235 14.535 ;
        RECT 177.150 13.495 177.530 13.875 ;
        RECT 178.935 13.495 179.315 13.875 ;
        RECT 181.790 13.495 182.170 13.875 ;
        RECT 183.575 13.495 183.955 13.875 ;
        RECT 186.430 13.495 186.810 13.875 ;
        RECT 188.215 13.495 188.595 13.875 ;
        RECT 191.070 13.495 191.450 13.875 ;
        RECT 192.855 13.495 193.235 13.875 ;
        RECT 177.150 12.835 177.530 13.215 ;
        RECT 178.935 12.835 179.315 13.215 ;
        RECT 181.790 12.835 182.170 13.215 ;
        RECT 183.575 12.835 183.955 13.215 ;
        RECT 186.430 12.835 186.810 13.215 ;
        RECT 188.215 12.835 188.595 13.215 ;
        RECT 191.070 12.835 191.450 13.215 ;
        RECT 192.855 12.835 193.235 13.215 ;
        RECT 177.150 12.175 177.530 12.555 ;
        RECT 178.935 12.175 179.315 12.555 ;
        RECT 181.790 12.175 182.170 12.555 ;
        RECT 183.575 12.175 183.955 12.555 ;
        RECT 186.430 12.175 186.810 12.555 ;
        RECT 188.215 12.175 188.595 12.555 ;
        RECT 191.070 12.175 191.450 12.555 ;
        RECT 192.855 12.175 193.235 12.555 ;
        RECT 177.150 11.515 177.530 11.895 ;
        RECT 178.935 11.515 179.315 11.895 ;
        RECT 181.790 11.515 182.170 11.895 ;
        RECT 183.575 11.515 183.955 11.895 ;
        RECT 186.430 11.515 186.810 11.895 ;
        RECT 188.215 11.515 188.595 11.895 ;
        RECT 191.070 11.515 191.450 11.895 ;
        RECT 192.855 11.515 193.235 11.895 ;
        RECT 177.150 10.855 177.530 11.235 ;
        RECT 178.935 10.855 179.315 11.235 ;
        RECT 181.790 10.855 182.170 11.235 ;
        RECT 183.575 10.855 183.955 11.235 ;
        RECT 186.430 10.855 186.810 11.235 ;
        RECT 188.215 10.855 188.595 11.235 ;
        RECT 191.070 10.855 191.450 11.235 ;
        RECT 192.855 10.855 193.235 11.235 ;
        RECT 177.150 10.195 177.530 10.575 ;
        RECT 178.935 10.195 179.315 10.575 ;
        RECT 181.790 10.195 182.170 10.575 ;
        RECT 183.575 10.195 183.955 10.575 ;
        RECT 186.430 10.195 186.810 10.575 ;
        RECT 188.215 10.195 188.595 10.575 ;
        RECT 191.070 10.195 191.450 10.575 ;
        RECT 192.855 10.195 193.235 10.575 ;
        RECT 177.150 9.535 177.530 9.915 ;
        RECT 178.935 9.535 179.315 9.915 ;
        RECT 181.790 9.535 182.170 9.915 ;
        RECT 183.575 9.535 183.955 9.915 ;
        RECT 186.430 9.535 186.810 9.915 ;
        RECT 188.215 9.535 188.595 9.915 ;
        RECT 191.070 9.535 191.450 9.915 ;
        RECT 192.855 9.535 193.235 9.915 ;
        RECT 177.150 8.875 177.530 9.255 ;
        RECT 178.935 8.875 179.315 9.255 ;
        RECT 181.790 8.875 182.170 9.255 ;
        RECT 183.575 8.875 183.955 9.255 ;
        RECT 186.430 8.875 186.810 9.255 ;
        RECT 188.215 8.875 188.595 9.255 ;
        RECT 191.070 8.875 191.450 9.255 ;
        RECT 192.855 8.875 193.235 9.255 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 42.110 8.090 42.490 8.470 ;
        RECT 56.940 8.090 57.320 8.470 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 42.110 7.430 42.490 7.810 ;
        RECT 56.940 7.430 57.320 7.810 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 42.110 6.770 42.490 7.150 ;
        RECT 56.940 6.770 57.320 7.150 ;
        RECT 0.850 4.690 1.230 5.070 ;
        RECT 1.990 4.690 2.370 5.070 ;
        RECT 8.030 4.720 8.410 5.100 ;
        RECT 8.690 4.720 9.070 5.100 ;
        RECT 9.350 4.720 9.730 5.100 ;
        RECT 14.560 4.690 14.940 5.070 ;
        RECT 15.220 4.690 15.600 5.070 ;
        RECT 15.880 4.690 16.260 5.070 ;
        RECT 17.920 4.690 18.300 5.070 ;
        RECT 18.580 4.690 18.960 5.070 ;
        RECT 19.240 4.690 19.620 5.070 ;
        RECT 26.220 4.720 26.600 5.100 ;
        RECT 26.880 4.720 27.260 5.100 ;
        RECT 27.540 4.720 27.920 5.100 ;
        RECT 32.750 4.690 33.130 5.070 ;
        RECT 33.410 4.690 33.790 5.070 ;
        RECT 34.070 4.690 34.450 5.070 ;
        RECT 36.110 4.690 36.490 5.070 ;
        RECT 36.770 4.690 37.150 5.070 ;
        RECT 37.430 4.690 37.810 5.070 ;
        RECT 39.490 4.690 39.870 5.070 ;
        RECT 45.530 4.720 45.910 5.100 ;
        RECT 46.190 4.720 46.570 5.100 ;
        RECT 46.850 4.720 47.230 5.100 ;
        RECT 52.060 4.690 52.440 5.070 ;
        RECT 52.720 4.690 53.100 5.070 ;
        RECT 53.380 4.690 53.760 5.070 ;
        RECT 60.360 4.720 60.740 5.100 ;
        RECT 61.020 4.720 61.400 5.100 ;
        RECT 61.680 4.720 62.060 5.100 ;
        RECT 66.890 4.690 67.270 5.070 ;
        RECT 67.550 4.690 67.930 5.070 ;
        RECT 68.210 4.690 68.590 5.070 ;
        RECT 70.250 4.690 70.630 5.070 ;
        RECT 70.910 4.690 71.290 5.070 ;
        RECT 71.570 4.690 71.950 5.070 ;
        RECT 73.630 4.690 74.010 5.070 ;
        RECT 74.630 4.690 75.010 5.070 ;
        RECT 75.290 4.690 75.670 5.070 ;
        RECT 75.950 4.690 76.330 5.070 ;
        RECT 76.870 4.690 77.250 5.070 ;
        RECT 77.530 4.690 77.910 5.070 ;
        RECT 78.190 4.690 78.570 5.070 ;
        RECT 79.210 4.690 79.590 5.070 ;
        RECT 79.870 4.690 80.250 5.070 ;
        RECT 80.530 4.690 80.910 5.070 ;
        RECT 82.470 4.690 82.850 5.070 ;
        RECT 83.130 4.690 83.510 5.070 ;
        RECT 83.790 4.690 84.170 5.070 ;
        RECT 84.710 4.690 85.090 5.070 ;
        RECT 85.370 4.690 85.750 5.070 ;
        RECT 86.030 4.690 86.410 5.070 ;
        RECT 86.950 4.690 87.330 5.070 ;
        RECT 87.610 4.690 87.990 5.070 ;
        RECT 88.270 4.690 88.650 5.070 ;
        RECT 89.190 4.690 89.570 5.070 ;
        RECT 89.850 4.690 90.230 5.070 ;
        RECT 90.510 4.690 90.890 5.070 ;
        RECT 91.430 4.690 91.810 5.070 ;
        RECT 92.090 4.690 92.470 5.070 ;
        RECT 92.750 4.690 93.130 5.070 ;
        RECT 93.790 4.690 94.170 5.070 ;
        RECT 94.790 4.690 95.170 5.070 ;
        RECT 95.450 4.690 95.830 5.070 ;
        RECT 96.110 4.690 96.490 5.070 ;
        RECT 97.030 4.690 97.410 5.070 ;
        RECT 97.690 4.690 98.070 5.070 ;
        RECT 98.350 4.690 98.730 5.070 ;
        RECT 99.270 4.690 99.650 5.070 ;
        RECT 99.930 4.690 100.310 5.070 ;
        RECT 100.590 4.690 100.970 5.070 ;
        RECT 101.610 4.690 101.990 5.070 ;
        RECT 102.270 4.690 102.650 5.070 ;
        RECT 102.930 4.690 103.310 5.070 ;
        RECT 104.870 4.690 105.250 5.070 ;
        RECT 105.530 4.690 105.910 5.070 ;
        RECT 106.190 4.690 106.570 5.070 ;
        RECT 107.110 4.690 107.490 5.070 ;
        RECT 107.770 4.690 108.150 5.070 ;
        RECT 108.430 4.690 108.810 5.070 ;
        RECT 109.350 4.690 109.730 5.070 ;
        RECT 110.010 4.690 110.390 5.070 ;
        RECT 110.670 4.690 111.050 5.070 ;
        RECT 111.590 4.690 111.970 5.070 ;
        RECT 112.250 4.690 112.630 5.070 ;
        RECT 112.910 4.690 113.290 5.070 ;
        RECT 113.950 4.690 114.330 5.070 ;
        RECT 114.950 4.690 115.330 5.070 ;
        RECT 115.610 4.690 115.990 5.070 ;
        RECT 116.270 4.690 116.650 5.070 ;
        RECT 117.190 4.690 117.570 5.070 ;
        RECT 117.850 4.690 118.230 5.070 ;
        RECT 118.510 4.690 118.890 5.070 ;
        RECT 119.430 4.690 119.810 5.070 ;
        RECT 120.090 4.690 120.470 5.070 ;
        RECT 120.750 4.690 121.130 5.070 ;
        RECT 121.770 4.690 122.150 5.070 ;
        RECT 122.430 4.690 122.810 5.070 ;
        RECT 123.090 4.690 123.470 5.070 ;
        RECT 125.030 4.690 125.410 5.070 ;
        RECT 125.690 4.690 126.070 5.070 ;
        RECT 126.350 4.690 126.730 5.070 ;
        RECT 127.270 4.690 127.650 5.070 ;
        RECT 127.930 4.690 128.310 5.070 ;
        RECT 128.590 4.690 128.970 5.070 ;
        RECT 129.510 4.690 129.890 5.070 ;
        RECT 130.170 4.690 130.550 5.070 ;
        RECT 130.830 4.690 131.210 5.070 ;
        RECT 131.750 4.690 132.130 5.070 ;
        RECT 132.410 4.690 132.790 5.070 ;
        RECT 133.070 4.690 133.450 5.070 ;
        RECT 134.110 4.690 134.490 5.070 ;
        RECT 135.110 4.690 135.490 5.070 ;
        RECT 135.770 4.690 136.150 5.070 ;
        RECT 136.430 4.690 136.810 5.070 ;
        RECT 137.350 4.690 137.730 5.070 ;
        RECT 138.010 4.690 138.390 5.070 ;
        RECT 138.670 4.690 139.050 5.070 ;
        RECT 139.590 4.690 139.970 5.070 ;
        RECT 140.250 4.690 140.630 5.070 ;
        RECT 140.910 4.690 141.290 5.070 ;
        RECT 141.830 4.690 142.210 5.070 ;
        RECT 142.490 4.690 142.870 5.070 ;
        RECT 143.150 4.690 143.530 5.070 ;
        RECT 144.170 4.690 144.550 5.070 ;
        RECT 144.830 4.690 145.210 5.070 ;
        RECT 145.490 4.690 145.870 5.070 ;
        RECT 147.430 4.690 147.810 5.070 ;
        RECT 148.090 4.690 148.470 5.070 ;
        RECT 148.750 4.690 149.130 5.070 ;
        RECT 149.670 4.690 150.050 5.070 ;
        RECT 150.330 4.690 150.710 5.070 ;
        RECT 150.990 4.690 151.370 5.070 ;
        RECT 151.910 4.690 152.290 5.070 ;
        RECT 152.570 4.690 152.950 5.070 ;
        RECT 153.230 4.690 153.610 5.070 ;
        RECT 154.270 4.690 154.650 5.070 ;
        RECT 155.270 4.690 155.650 5.070 ;
        RECT 155.930 4.690 156.310 5.070 ;
        RECT 156.590 4.690 156.970 5.070 ;
        RECT 157.510 4.690 157.890 5.070 ;
        RECT 158.170 4.690 158.550 5.070 ;
        RECT 158.830 4.690 159.210 5.070 ;
        RECT 159.750 4.690 160.130 5.070 ;
        RECT 160.410 4.690 160.790 5.070 ;
        RECT 161.070 4.690 161.450 5.070 ;
        RECT 161.990 4.690 162.370 5.070 ;
        RECT 162.650 4.690 163.030 5.070 ;
        RECT 163.310 4.690 163.690 5.070 ;
        RECT 164.230 4.690 164.610 5.070 ;
        RECT 164.890 4.690 165.270 5.070 ;
        RECT 165.550 4.690 165.930 5.070 ;
        RECT 166.570 4.690 166.950 5.070 ;
        RECT 167.230 4.690 167.610 5.070 ;
        RECT 167.890 4.690 168.270 5.070 ;
        RECT 169.830 4.690 170.210 5.070 ;
        RECT 170.490 4.690 170.870 5.070 ;
        RECT 171.150 4.690 171.530 5.070 ;
        RECT 172.070 4.690 172.450 5.070 ;
        RECT 172.730 4.690 173.110 5.070 ;
        RECT 173.390 4.690 173.770 5.070 ;
        RECT 174.410 4.690 174.790 5.070 ;
        RECT 0.850 0.770 1.230 1.150 ;
        RECT 1.990 0.770 2.370 1.150 ;
        RECT 7.430 0.770 7.810 1.150 ;
        RECT 8.090 0.770 8.470 1.150 ;
        RECT 8.750 0.770 9.130 1.150 ;
        RECT 14.300 0.770 14.680 1.150 ;
        RECT 15.620 0.770 16.000 1.150 ;
        RECT 17.660 0.770 18.040 1.150 ;
        RECT 18.980 0.770 19.360 1.150 ;
        RECT 25.620 0.770 26.000 1.150 ;
        RECT 26.280 0.770 26.660 1.150 ;
        RECT 26.940 0.770 27.320 1.150 ;
        RECT 32.490 0.770 32.870 1.150 ;
        RECT 33.810 0.770 34.190 1.150 ;
        RECT 35.850 0.770 36.230 1.150 ;
        RECT 37.170 0.770 37.550 1.150 ;
        RECT 39.490 0.770 39.870 1.150 ;
        RECT 44.930 0.770 45.310 1.150 ;
        RECT 45.590 0.770 45.970 1.150 ;
        RECT 46.250 0.770 46.630 1.150 ;
        RECT 51.800 0.770 52.180 1.150 ;
        RECT 53.120 0.770 53.500 1.150 ;
        RECT 59.760 0.770 60.140 1.150 ;
        RECT 60.420 0.770 60.800 1.150 ;
        RECT 61.080 0.770 61.460 1.150 ;
        RECT 66.630 0.770 67.010 1.150 ;
        RECT 67.950 0.770 68.330 1.150 ;
        RECT 69.990 0.770 70.370 1.150 ;
        RECT 71.310 0.770 71.690 1.150 ;
        RECT 73.630 0.770 74.010 1.150 ;
        RECT 74.630 0.770 75.010 1.150 ;
        RECT 75.290 0.770 75.670 1.150 ;
        RECT 75.950 0.770 76.330 1.150 ;
        RECT 76.870 0.770 77.250 1.150 ;
        RECT 77.530 0.770 77.910 1.150 ;
        RECT 78.190 0.770 78.570 1.150 ;
        RECT 78.950 0.770 79.330 1.150 ;
        RECT 80.270 0.770 80.650 1.150 ;
        RECT 82.470 0.770 82.850 1.150 ;
        RECT 83.130 0.770 83.510 1.150 ;
        RECT 83.790 0.770 84.170 1.150 ;
        RECT 84.710 0.770 85.090 1.150 ;
        RECT 85.370 0.770 85.750 1.150 ;
        RECT 86.030 0.770 86.410 1.150 ;
        RECT 86.950 0.770 87.330 1.150 ;
        RECT 87.610 0.770 87.990 1.150 ;
        RECT 88.270 0.770 88.650 1.150 ;
        RECT 89.190 0.770 89.570 1.150 ;
        RECT 89.850 0.770 90.230 1.150 ;
        RECT 90.510 0.770 90.890 1.150 ;
        RECT 91.430 0.770 91.810 1.150 ;
        RECT 92.090 0.770 92.470 1.150 ;
        RECT 92.750 0.770 93.130 1.150 ;
        RECT 93.790 0.770 94.170 1.150 ;
        RECT 94.790 0.770 95.170 1.150 ;
        RECT 95.450 0.770 95.830 1.150 ;
        RECT 96.110 0.770 96.490 1.150 ;
        RECT 97.030 0.770 97.410 1.150 ;
        RECT 97.690 0.770 98.070 1.150 ;
        RECT 98.350 0.770 98.730 1.150 ;
        RECT 99.270 0.770 99.650 1.150 ;
        RECT 99.930 0.770 100.310 1.150 ;
        RECT 100.590 0.770 100.970 1.150 ;
        RECT 101.350 0.770 101.730 1.150 ;
        RECT 102.670 0.770 103.050 1.150 ;
        RECT 104.870 0.770 105.250 1.150 ;
        RECT 105.530 0.770 105.910 1.150 ;
        RECT 106.190 0.770 106.570 1.150 ;
        RECT 107.110 0.770 107.490 1.150 ;
        RECT 107.770 0.770 108.150 1.150 ;
        RECT 108.430 0.770 108.810 1.150 ;
        RECT 109.350 0.770 109.730 1.150 ;
        RECT 110.010 0.770 110.390 1.150 ;
        RECT 110.670 0.770 111.050 1.150 ;
        RECT 111.590 0.770 111.970 1.150 ;
        RECT 112.250 0.770 112.630 1.150 ;
        RECT 112.910 0.770 113.290 1.150 ;
        RECT 113.950 0.770 114.330 1.150 ;
        RECT 114.950 0.770 115.330 1.150 ;
        RECT 115.610 0.770 115.990 1.150 ;
        RECT 116.270 0.770 116.650 1.150 ;
        RECT 117.190 0.770 117.570 1.150 ;
        RECT 117.850 0.770 118.230 1.150 ;
        RECT 118.510 0.770 118.890 1.150 ;
        RECT 119.430 0.770 119.810 1.150 ;
        RECT 120.090 0.770 120.470 1.150 ;
        RECT 120.750 0.770 121.130 1.150 ;
        RECT 121.510 0.770 121.890 1.150 ;
        RECT 122.830 0.770 123.210 1.150 ;
        RECT 125.030 0.770 125.410 1.150 ;
        RECT 125.690 0.770 126.070 1.150 ;
        RECT 126.350 0.770 126.730 1.150 ;
        RECT 127.270 0.770 127.650 1.150 ;
        RECT 127.930 0.770 128.310 1.150 ;
        RECT 128.590 0.770 128.970 1.150 ;
        RECT 129.510 0.770 129.890 1.150 ;
        RECT 130.170 0.770 130.550 1.150 ;
        RECT 130.830 0.770 131.210 1.150 ;
        RECT 131.750 0.770 132.130 1.150 ;
        RECT 132.410 0.770 132.790 1.150 ;
        RECT 133.070 0.770 133.450 1.150 ;
        RECT 134.110 0.770 134.490 1.150 ;
        RECT 135.110 0.770 135.490 1.150 ;
        RECT 135.770 0.770 136.150 1.150 ;
        RECT 136.430 0.770 136.810 1.150 ;
        RECT 137.350 0.770 137.730 1.150 ;
        RECT 138.010 0.770 138.390 1.150 ;
        RECT 138.670 0.770 139.050 1.150 ;
        RECT 139.590 0.770 139.970 1.150 ;
        RECT 140.250 0.770 140.630 1.150 ;
        RECT 140.910 0.770 141.290 1.150 ;
        RECT 141.830 0.770 142.210 1.150 ;
        RECT 142.490 0.770 142.870 1.150 ;
        RECT 143.150 0.770 143.530 1.150 ;
        RECT 143.910 0.770 144.290 1.150 ;
        RECT 145.230 0.770 145.610 1.150 ;
        RECT 147.430 0.770 147.810 1.150 ;
        RECT 148.090 0.770 148.470 1.150 ;
        RECT 148.750 0.770 149.130 1.150 ;
        RECT 149.670 0.770 150.050 1.150 ;
        RECT 150.330 0.770 150.710 1.150 ;
        RECT 150.990 0.770 151.370 1.150 ;
        RECT 151.910 0.770 152.290 1.150 ;
        RECT 152.570 0.770 152.950 1.150 ;
        RECT 153.230 0.770 153.610 1.150 ;
        RECT 154.270 0.770 154.650 1.150 ;
        RECT 155.270 0.770 155.650 1.150 ;
        RECT 155.930 0.770 156.310 1.150 ;
        RECT 156.590 0.770 156.970 1.150 ;
        RECT 157.510 0.770 157.890 1.150 ;
        RECT 158.170 0.770 158.550 1.150 ;
        RECT 158.830 0.770 159.210 1.150 ;
        RECT 159.750 0.770 160.130 1.150 ;
        RECT 160.410 0.770 160.790 1.150 ;
        RECT 161.070 0.770 161.450 1.150 ;
        RECT 161.990 0.770 162.370 1.150 ;
        RECT 162.650 0.770 163.030 1.150 ;
        RECT 163.310 0.770 163.690 1.150 ;
        RECT 164.230 0.770 164.610 1.150 ;
        RECT 164.890 0.770 165.270 1.150 ;
        RECT 165.550 0.770 165.930 1.150 ;
        RECT 166.310 0.770 166.690 1.150 ;
        RECT 167.630 0.770 168.010 1.150 ;
        RECT 169.830 0.770 170.210 1.150 ;
        RECT 170.490 0.770 170.870 1.150 ;
        RECT 171.150 0.770 171.530 1.150 ;
        RECT 172.070 0.770 172.450 1.150 ;
        RECT 172.730 0.770 173.110 1.150 ;
        RECT 173.390 0.770 173.770 1.150 ;
        RECT 174.410 0.770 174.790 1.150 ;
      LAYER Via3 ;
        RECT 0.815 58.795 1.095 59.075 ;
        RECT 11.105 58.795 11.385 59.075 ;
        RECT 21.390 58.795 21.670 59.075 ;
        RECT 22.810 58.795 23.090 59.075 ;
        RECT 33.100 58.795 33.380 59.075 ;
        RECT 43.385 58.795 43.665 59.075 ;
        RECT 44.805 58.795 45.085 59.075 ;
        RECT 55.095 58.795 55.375 59.075 ;
        RECT 65.380 58.795 65.660 59.075 ;
        RECT 66.800 58.795 67.080 59.075 ;
        RECT 77.090 58.795 77.370 59.075 ;
        RECT 87.375 58.795 87.655 59.075 ;
        RECT 88.795 58.795 89.075 59.075 ;
        RECT 99.085 58.795 99.365 59.075 ;
        RECT 109.370 58.795 109.650 59.075 ;
        RECT 110.790 58.795 111.070 59.075 ;
        RECT 121.080 58.795 121.360 59.075 ;
        RECT 131.365 58.795 131.645 59.075 ;
        RECT 132.785 58.795 133.065 59.075 ;
        RECT 143.075 58.795 143.355 59.075 ;
        RECT 153.360 58.795 153.640 59.075 ;
        RECT 154.780 58.795 155.060 59.075 ;
        RECT 165.070 58.795 165.350 59.075 ;
        RECT 175.355 58.795 175.635 59.075 ;
        RECT 0.815 58.135 1.095 58.415 ;
        RECT 11.105 58.135 11.385 58.415 ;
        RECT 21.390 58.135 21.670 58.415 ;
        RECT 22.810 58.135 23.090 58.415 ;
        RECT 33.100 58.135 33.380 58.415 ;
        RECT 43.385 58.135 43.665 58.415 ;
        RECT 44.805 58.135 45.085 58.415 ;
        RECT 55.095 58.135 55.375 58.415 ;
        RECT 65.380 58.135 65.660 58.415 ;
        RECT 66.800 58.135 67.080 58.415 ;
        RECT 77.090 58.135 77.370 58.415 ;
        RECT 87.375 58.135 87.655 58.415 ;
        RECT 88.795 58.135 89.075 58.415 ;
        RECT 99.085 58.135 99.365 58.415 ;
        RECT 109.370 58.135 109.650 58.415 ;
        RECT 110.790 58.135 111.070 58.415 ;
        RECT 121.080 58.135 121.360 58.415 ;
        RECT 131.365 58.135 131.645 58.415 ;
        RECT 132.785 58.135 133.065 58.415 ;
        RECT 143.075 58.135 143.355 58.415 ;
        RECT 153.360 58.135 153.640 58.415 ;
        RECT 154.780 58.135 155.060 58.415 ;
        RECT 165.070 58.135 165.350 58.415 ;
        RECT 175.355 58.135 175.635 58.415 ;
        RECT 0.815 57.475 1.095 57.755 ;
        RECT 11.105 57.475 11.385 57.755 ;
        RECT 21.390 57.475 21.670 57.755 ;
        RECT 22.810 57.475 23.090 57.755 ;
        RECT 33.100 57.475 33.380 57.755 ;
        RECT 43.385 57.475 43.665 57.755 ;
        RECT 44.805 57.475 45.085 57.755 ;
        RECT 55.095 57.475 55.375 57.755 ;
        RECT 65.380 57.475 65.660 57.755 ;
        RECT 66.800 57.475 67.080 57.755 ;
        RECT 77.090 57.475 77.370 57.755 ;
        RECT 87.375 57.475 87.655 57.755 ;
        RECT 88.795 57.475 89.075 57.755 ;
        RECT 99.085 57.475 99.365 57.755 ;
        RECT 109.370 57.475 109.650 57.755 ;
        RECT 110.790 57.475 111.070 57.755 ;
        RECT 121.080 57.475 121.360 57.755 ;
        RECT 131.365 57.475 131.645 57.755 ;
        RECT 132.785 57.475 133.065 57.755 ;
        RECT 143.075 57.475 143.355 57.755 ;
        RECT 153.360 57.475 153.640 57.755 ;
        RECT 154.780 57.475 155.060 57.755 ;
        RECT 165.070 57.475 165.350 57.755 ;
        RECT 175.355 57.475 175.635 57.755 ;
        RECT 0.815 56.815 1.095 57.095 ;
        RECT 11.105 56.815 11.385 57.095 ;
        RECT 21.390 56.815 21.670 57.095 ;
        RECT 22.810 56.815 23.090 57.095 ;
        RECT 33.100 56.815 33.380 57.095 ;
        RECT 43.385 56.815 43.665 57.095 ;
        RECT 44.805 56.815 45.085 57.095 ;
        RECT 55.095 56.815 55.375 57.095 ;
        RECT 65.380 56.815 65.660 57.095 ;
        RECT 66.800 56.815 67.080 57.095 ;
        RECT 77.090 56.815 77.370 57.095 ;
        RECT 87.375 56.815 87.655 57.095 ;
        RECT 88.795 56.815 89.075 57.095 ;
        RECT 99.085 56.815 99.365 57.095 ;
        RECT 109.370 56.815 109.650 57.095 ;
        RECT 110.790 56.815 111.070 57.095 ;
        RECT 121.080 56.815 121.360 57.095 ;
        RECT 131.365 56.815 131.645 57.095 ;
        RECT 132.785 56.815 133.065 57.095 ;
        RECT 143.075 56.815 143.355 57.095 ;
        RECT 153.360 56.815 153.640 57.095 ;
        RECT 154.780 56.815 155.060 57.095 ;
        RECT 165.070 56.815 165.350 57.095 ;
        RECT 175.355 56.815 175.635 57.095 ;
        RECT 0.815 56.155 1.095 56.435 ;
        RECT 11.105 56.155 11.385 56.435 ;
        RECT 21.390 56.155 21.670 56.435 ;
        RECT 22.810 56.155 23.090 56.435 ;
        RECT 33.100 56.155 33.380 56.435 ;
        RECT 43.385 56.155 43.665 56.435 ;
        RECT 44.805 56.155 45.085 56.435 ;
        RECT 55.095 56.155 55.375 56.435 ;
        RECT 65.380 56.155 65.660 56.435 ;
        RECT 66.800 56.155 67.080 56.435 ;
        RECT 77.090 56.155 77.370 56.435 ;
        RECT 87.375 56.155 87.655 56.435 ;
        RECT 88.795 56.155 89.075 56.435 ;
        RECT 99.085 56.155 99.365 56.435 ;
        RECT 109.370 56.155 109.650 56.435 ;
        RECT 110.790 56.155 111.070 56.435 ;
        RECT 121.080 56.155 121.360 56.435 ;
        RECT 131.365 56.155 131.645 56.435 ;
        RECT 132.785 56.155 133.065 56.435 ;
        RECT 143.075 56.155 143.355 56.435 ;
        RECT 153.360 56.155 153.640 56.435 ;
        RECT 154.780 56.155 155.060 56.435 ;
        RECT 165.070 56.155 165.350 56.435 ;
        RECT 175.355 56.155 175.635 56.435 ;
        RECT 0.815 55.495 1.095 55.775 ;
        RECT 11.105 55.495 11.385 55.775 ;
        RECT 21.390 55.495 21.670 55.775 ;
        RECT 22.810 55.495 23.090 55.775 ;
        RECT 33.100 55.495 33.380 55.775 ;
        RECT 43.385 55.495 43.665 55.775 ;
        RECT 44.805 55.495 45.085 55.775 ;
        RECT 55.095 55.495 55.375 55.775 ;
        RECT 65.380 55.495 65.660 55.775 ;
        RECT 66.800 55.495 67.080 55.775 ;
        RECT 77.090 55.495 77.370 55.775 ;
        RECT 87.375 55.495 87.655 55.775 ;
        RECT 88.795 55.495 89.075 55.775 ;
        RECT 99.085 55.495 99.365 55.775 ;
        RECT 109.370 55.495 109.650 55.775 ;
        RECT 110.790 55.495 111.070 55.775 ;
        RECT 121.080 55.495 121.360 55.775 ;
        RECT 131.365 55.495 131.645 55.775 ;
        RECT 132.785 55.495 133.065 55.775 ;
        RECT 143.075 55.495 143.355 55.775 ;
        RECT 153.360 55.495 153.640 55.775 ;
        RECT 154.780 55.495 155.060 55.775 ;
        RECT 165.070 55.495 165.350 55.775 ;
        RECT 175.355 55.495 175.635 55.775 ;
        RECT 177.200 55.165 177.480 55.445 ;
        RECT 0.815 54.835 1.095 55.115 ;
        RECT 11.105 54.835 11.385 55.115 ;
        RECT 21.390 54.835 21.670 55.115 ;
        RECT 22.810 54.835 23.090 55.115 ;
        RECT 33.100 54.835 33.380 55.115 ;
        RECT 43.385 54.835 43.665 55.115 ;
        RECT 44.805 54.835 45.085 55.115 ;
        RECT 55.095 54.835 55.375 55.115 ;
        RECT 65.380 54.835 65.660 55.115 ;
        RECT 66.800 54.835 67.080 55.115 ;
        RECT 77.090 54.835 77.370 55.115 ;
        RECT 87.375 54.835 87.655 55.115 ;
        RECT 88.795 54.835 89.075 55.115 ;
        RECT 99.085 54.835 99.365 55.115 ;
        RECT 109.370 54.835 109.650 55.115 ;
        RECT 110.790 54.835 111.070 55.115 ;
        RECT 121.080 54.835 121.360 55.115 ;
        RECT 131.365 54.835 131.645 55.115 ;
        RECT 132.785 54.835 133.065 55.115 ;
        RECT 143.075 54.835 143.355 55.115 ;
        RECT 153.360 54.835 153.640 55.115 ;
        RECT 154.780 54.835 155.060 55.115 ;
        RECT 165.070 54.835 165.350 55.115 ;
        RECT 178.985 55.165 179.265 55.445 ;
        RECT 181.840 55.165 182.120 55.445 ;
        RECT 183.625 55.165 183.905 55.445 ;
        RECT 186.480 55.165 186.760 55.445 ;
        RECT 188.265 55.165 188.545 55.445 ;
        RECT 191.120 55.165 191.400 55.445 ;
        RECT 192.905 55.165 193.185 55.445 ;
        RECT 175.355 54.835 175.635 55.115 ;
        RECT 177.200 54.505 177.480 54.785 ;
        RECT 0.815 54.175 1.095 54.455 ;
        RECT 11.105 54.175 11.385 54.455 ;
        RECT 21.390 54.175 21.670 54.455 ;
        RECT 22.810 54.175 23.090 54.455 ;
        RECT 33.100 54.175 33.380 54.455 ;
        RECT 43.385 54.175 43.665 54.455 ;
        RECT 44.805 54.175 45.085 54.455 ;
        RECT 55.095 54.175 55.375 54.455 ;
        RECT 65.380 54.175 65.660 54.455 ;
        RECT 66.800 54.175 67.080 54.455 ;
        RECT 77.090 54.175 77.370 54.455 ;
        RECT 87.375 54.175 87.655 54.455 ;
        RECT 88.795 54.175 89.075 54.455 ;
        RECT 99.085 54.175 99.365 54.455 ;
        RECT 109.370 54.175 109.650 54.455 ;
        RECT 110.790 54.175 111.070 54.455 ;
        RECT 121.080 54.175 121.360 54.455 ;
        RECT 131.365 54.175 131.645 54.455 ;
        RECT 132.785 54.175 133.065 54.455 ;
        RECT 143.075 54.175 143.355 54.455 ;
        RECT 153.360 54.175 153.640 54.455 ;
        RECT 154.780 54.175 155.060 54.455 ;
        RECT 165.070 54.175 165.350 54.455 ;
        RECT 178.985 54.505 179.265 54.785 ;
        RECT 181.840 54.505 182.120 54.785 ;
        RECT 183.625 54.505 183.905 54.785 ;
        RECT 186.480 54.505 186.760 54.785 ;
        RECT 188.265 54.505 188.545 54.785 ;
        RECT 191.120 54.505 191.400 54.785 ;
        RECT 192.905 54.505 193.185 54.785 ;
        RECT 175.355 54.175 175.635 54.455 ;
        RECT 177.200 53.845 177.480 54.125 ;
        RECT 0.815 53.515 1.095 53.795 ;
        RECT 11.105 53.515 11.385 53.795 ;
        RECT 21.390 53.515 21.670 53.795 ;
        RECT 22.810 53.515 23.090 53.795 ;
        RECT 33.100 53.515 33.380 53.795 ;
        RECT 43.385 53.515 43.665 53.795 ;
        RECT 44.805 53.515 45.085 53.795 ;
        RECT 55.095 53.515 55.375 53.795 ;
        RECT 65.380 53.515 65.660 53.795 ;
        RECT 66.800 53.515 67.080 53.795 ;
        RECT 77.090 53.515 77.370 53.795 ;
        RECT 87.375 53.515 87.655 53.795 ;
        RECT 88.795 53.515 89.075 53.795 ;
        RECT 99.085 53.515 99.365 53.795 ;
        RECT 109.370 53.515 109.650 53.795 ;
        RECT 110.790 53.515 111.070 53.795 ;
        RECT 121.080 53.515 121.360 53.795 ;
        RECT 131.365 53.515 131.645 53.795 ;
        RECT 132.785 53.515 133.065 53.795 ;
        RECT 143.075 53.515 143.355 53.795 ;
        RECT 153.360 53.515 153.640 53.795 ;
        RECT 154.780 53.515 155.060 53.795 ;
        RECT 165.070 53.515 165.350 53.795 ;
        RECT 178.985 53.845 179.265 54.125 ;
        RECT 181.840 53.845 182.120 54.125 ;
        RECT 183.625 53.845 183.905 54.125 ;
        RECT 186.480 53.845 186.760 54.125 ;
        RECT 188.265 53.845 188.545 54.125 ;
        RECT 191.120 53.845 191.400 54.125 ;
        RECT 192.905 53.845 193.185 54.125 ;
        RECT 175.355 53.515 175.635 53.795 ;
        RECT 177.200 53.185 177.480 53.465 ;
        RECT 0.815 52.855 1.095 53.135 ;
        RECT 11.105 52.855 11.385 53.135 ;
        RECT 21.390 52.855 21.670 53.135 ;
        RECT 22.810 52.855 23.090 53.135 ;
        RECT 33.100 52.855 33.380 53.135 ;
        RECT 43.385 52.855 43.665 53.135 ;
        RECT 44.805 52.855 45.085 53.135 ;
        RECT 55.095 52.855 55.375 53.135 ;
        RECT 65.380 52.855 65.660 53.135 ;
        RECT 66.800 52.855 67.080 53.135 ;
        RECT 77.090 52.855 77.370 53.135 ;
        RECT 87.375 52.855 87.655 53.135 ;
        RECT 88.795 52.855 89.075 53.135 ;
        RECT 99.085 52.855 99.365 53.135 ;
        RECT 109.370 52.855 109.650 53.135 ;
        RECT 110.790 52.855 111.070 53.135 ;
        RECT 121.080 52.855 121.360 53.135 ;
        RECT 131.365 52.855 131.645 53.135 ;
        RECT 132.785 52.855 133.065 53.135 ;
        RECT 143.075 52.855 143.355 53.135 ;
        RECT 153.360 52.855 153.640 53.135 ;
        RECT 154.780 52.855 155.060 53.135 ;
        RECT 165.070 52.855 165.350 53.135 ;
        RECT 178.985 53.185 179.265 53.465 ;
        RECT 181.840 53.185 182.120 53.465 ;
        RECT 183.625 53.185 183.905 53.465 ;
        RECT 186.480 53.185 186.760 53.465 ;
        RECT 188.265 53.185 188.545 53.465 ;
        RECT 191.120 53.185 191.400 53.465 ;
        RECT 192.905 53.185 193.185 53.465 ;
        RECT 175.355 52.855 175.635 53.135 ;
        RECT 177.200 52.525 177.480 52.805 ;
        RECT 0.815 52.195 1.095 52.475 ;
        RECT 11.105 52.195 11.385 52.475 ;
        RECT 21.390 52.195 21.670 52.475 ;
        RECT 22.810 52.195 23.090 52.475 ;
        RECT 33.100 52.195 33.380 52.475 ;
        RECT 43.385 52.195 43.665 52.475 ;
        RECT 44.805 52.195 45.085 52.475 ;
        RECT 55.095 52.195 55.375 52.475 ;
        RECT 65.380 52.195 65.660 52.475 ;
        RECT 66.800 52.195 67.080 52.475 ;
        RECT 77.090 52.195 77.370 52.475 ;
        RECT 87.375 52.195 87.655 52.475 ;
        RECT 88.795 52.195 89.075 52.475 ;
        RECT 99.085 52.195 99.365 52.475 ;
        RECT 109.370 52.195 109.650 52.475 ;
        RECT 110.790 52.195 111.070 52.475 ;
        RECT 121.080 52.195 121.360 52.475 ;
        RECT 131.365 52.195 131.645 52.475 ;
        RECT 132.785 52.195 133.065 52.475 ;
        RECT 143.075 52.195 143.355 52.475 ;
        RECT 153.360 52.195 153.640 52.475 ;
        RECT 154.780 52.195 155.060 52.475 ;
        RECT 165.070 52.195 165.350 52.475 ;
        RECT 178.985 52.525 179.265 52.805 ;
        RECT 181.840 52.525 182.120 52.805 ;
        RECT 183.625 52.525 183.905 52.805 ;
        RECT 186.480 52.525 186.760 52.805 ;
        RECT 188.265 52.525 188.545 52.805 ;
        RECT 191.120 52.525 191.400 52.805 ;
        RECT 192.905 52.525 193.185 52.805 ;
        RECT 175.355 52.195 175.635 52.475 ;
        RECT 177.200 51.865 177.480 52.145 ;
        RECT 0.815 51.535 1.095 51.815 ;
        RECT 11.105 51.535 11.385 51.815 ;
        RECT 21.390 51.535 21.670 51.815 ;
        RECT 22.810 51.535 23.090 51.815 ;
        RECT 33.100 51.535 33.380 51.815 ;
        RECT 43.385 51.535 43.665 51.815 ;
        RECT 44.805 51.535 45.085 51.815 ;
        RECT 55.095 51.535 55.375 51.815 ;
        RECT 65.380 51.535 65.660 51.815 ;
        RECT 66.800 51.535 67.080 51.815 ;
        RECT 77.090 51.535 77.370 51.815 ;
        RECT 87.375 51.535 87.655 51.815 ;
        RECT 88.795 51.535 89.075 51.815 ;
        RECT 99.085 51.535 99.365 51.815 ;
        RECT 109.370 51.535 109.650 51.815 ;
        RECT 110.790 51.535 111.070 51.815 ;
        RECT 121.080 51.535 121.360 51.815 ;
        RECT 131.365 51.535 131.645 51.815 ;
        RECT 132.785 51.535 133.065 51.815 ;
        RECT 143.075 51.535 143.355 51.815 ;
        RECT 153.360 51.535 153.640 51.815 ;
        RECT 154.780 51.535 155.060 51.815 ;
        RECT 165.070 51.535 165.350 51.815 ;
        RECT 178.985 51.865 179.265 52.145 ;
        RECT 181.840 51.865 182.120 52.145 ;
        RECT 183.625 51.865 183.905 52.145 ;
        RECT 186.480 51.865 186.760 52.145 ;
        RECT 188.265 51.865 188.545 52.145 ;
        RECT 191.120 51.865 191.400 52.145 ;
        RECT 192.905 51.865 193.185 52.145 ;
        RECT 175.355 51.535 175.635 51.815 ;
        RECT 177.200 51.205 177.480 51.485 ;
        RECT 0.815 50.875 1.095 51.155 ;
        RECT 11.105 50.875 11.385 51.155 ;
        RECT 21.390 50.875 21.670 51.155 ;
        RECT 22.810 50.875 23.090 51.155 ;
        RECT 33.100 50.875 33.380 51.155 ;
        RECT 43.385 50.875 43.665 51.155 ;
        RECT 44.805 50.875 45.085 51.155 ;
        RECT 55.095 50.875 55.375 51.155 ;
        RECT 65.380 50.875 65.660 51.155 ;
        RECT 66.800 50.875 67.080 51.155 ;
        RECT 77.090 50.875 77.370 51.155 ;
        RECT 87.375 50.875 87.655 51.155 ;
        RECT 88.795 50.875 89.075 51.155 ;
        RECT 99.085 50.875 99.365 51.155 ;
        RECT 109.370 50.875 109.650 51.155 ;
        RECT 110.790 50.875 111.070 51.155 ;
        RECT 121.080 50.875 121.360 51.155 ;
        RECT 131.365 50.875 131.645 51.155 ;
        RECT 132.785 50.875 133.065 51.155 ;
        RECT 143.075 50.875 143.355 51.155 ;
        RECT 153.360 50.875 153.640 51.155 ;
        RECT 154.780 50.875 155.060 51.155 ;
        RECT 165.070 50.875 165.350 51.155 ;
        RECT 178.985 51.205 179.265 51.485 ;
        RECT 181.840 51.205 182.120 51.485 ;
        RECT 183.625 51.205 183.905 51.485 ;
        RECT 186.480 51.205 186.760 51.485 ;
        RECT 188.265 51.205 188.545 51.485 ;
        RECT 191.120 51.205 191.400 51.485 ;
        RECT 192.905 51.205 193.185 51.485 ;
        RECT 175.355 50.875 175.635 51.155 ;
        RECT 177.200 50.545 177.480 50.825 ;
        RECT 0.815 50.215 1.095 50.495 ;
        RECT 11.105 50.215 11.385 50.495 ;
        RECT 21.390 50.215 21.670 50.495 ;
        RECT 22.810 50.215 23.090 50.495 ;
        RECT 33.100 50.215 33.380 50.495 ;
        RECT 43.385 50.215 43.665 50.495 ;
        RECT 44.805 50.215 45.085 50.495 ;
        RECT 55.095 50.215 55.375 50.495 ;
        RECT 65.380 50.215 65.660 50.495 ;
        RECT 66.800 50.215 67.080 50.495 ;
        RECT 77.090 50.215 77.370 50.495 ;
        RECT 87.375 50.215 87.655 50.495 ;
        RECT 88.795 50.215 89.075 50.495 ;
        RECT 99.085 50.215 99.365 50.495 ;
        RECT 109.370 50.215 109.650 50.495 ;
        RECT 110.790 50.215 111.070 50.495 ;
        RECT 121.080 50.215 121.360 50.495 ;
        RECT 131.365 50.215 131.645 50.495 ;
        RECT 132.785 50.215 133.065 50.495 ;
        RECT 143.075 50.215 143.355 50.495 ;
        RECT 153.360 50.215 153.640 50.495 ;
        RECT 154.780 50.215 155.060 50.495 ;
        RECT 165.070 50.215 165.350 50.495 ;
        RECT 178.985 50.545 179.265 50.825 ;
        RECT 181.840 50.545 182.120 50.825 ;
        RECT 183.625 50.545 183.905 50.825 ;
        RECT 186.480 50.545 186.760 50.825 ;
        RECT 188.265 50.545 188.545 50.825 ;
        RECT 191.120 50.545 191.400 50.825 ;
        RECT 192.905 50.545 193.185 50.825 ;
        RECT 175.355 50.215 175.635 50.495 ;
        RECT 4.660 47.855 4.940 48.135 ;
        RECT 4.660 47.195 4.940 47.475 ;
        RECT 4.660 46.535 4.940 46.815 ;
        RECT 56.990 45.155 57.270 45.435 ;
        RECT 56.990 44.495 57.270 44.775 ;
        RECT 56.990 43.835 57.270 44.115 ;
        RECT 42.160 24.955 42.440 25.235 ;
        RECT 42.160 24.295 42.440 24.575 ;
        RECT 42.160 23.635 42.440 23.915 ;
        RECT 22.850 22.255 23.130 22.535 ;
        RECT 22.850 21.595 23.130 21.875 ;
        RECT 22.850 20.935 23.130 21.215 ;
        RECT 177.200 18.165 177.480 18.445 ;
        RECT 178.985 18.165 179.265 18.445 ;
        RECT 181.840 18.165 182.120 18.445 ;
        RECT 183.625 18.165 183.905 18.445 ;
        RECT 186.480 18.165 186.760 18.445 ;
        RECT 188.265 18.165 188.545 18.445 ;
        RECT 191.120 18.165 191.400 18.445 ;
        RECT 192.905 18.165 193.185 18.445 ;
        RECT 177.200 17.505 177.480 17.785 ;
        RECT 178.985 17.505 179.265 17.785 ;
        RECT 181.840 17.505 182.120 17.785 ;
        RECT 183.625 17.505 183.905 17.785 ;
        RECT 186.480 17.505 186.760 17.785 ;
        RECT 188.265 17.505 188.545 17.785 ;
        RECT 191.120 17.505 191.400 17.785 ;
        RECT 192.905 17.505 193.185 17.785 ;
        RECT 177.200 16.845 177.480 17.125 ;
        RECT 178.985 16.845 179.265 17.125 ;
        RECT 181.840 16.845 182.120 17.125 ;
        RECT 183.625 16.845 183.905 17.125 ;
        RECT 186.480 16.845 186.760 17.125 ;
        RECT 188.265 16.845 188.545 17.125 ;
        RECT 191.120 16.845 191.400 17.125 ;
        RECT 192.905 16.845 193.185 17.125 ;
        RECT 177.200 16.185 177.480 16.465 ;
        RECT 178.985 16.185 179.265 16.465 ;
        RECT 181.840 16.185 182.120 16.465 ;
        RECT 183.625 16.185 183.905 16.465 ;
        RECT 186.480 16.185 186.760 16.465 ;
        RECT 188.265 16.185 188.545 16.465 ;
        RECT 191.120 16.185 191.400 16.465 ;
        RECT 192.905 16.185 193.185 16.465 ;
        RECT 177.200 15.525 177.480 15.805 ;
        RECT 178.985 15.525 179.265 15.805 ;
        RECT 181.840 15.525 182.120 15.805 ;
        RECT 183.625 15.525 183.905 15.805 ;
        RECT 186.480 15.525 186.760 15.805 ;
        RECT 188.265 15.525 188.545 15.805 ;
        RECT 191.120 15.525 191.400 15.805 ;
        RECT 192.905 15.525 193.185 15.805 ;
        RECT 177.200 14.865 177.480 15.145 ;
        RECT 178.985 14.865 179.265 15.145 ;
        RECT 181.840 14.865 182.120 15.145 ;
        RECT 183.625 14.865 183.905 15.145 ;
        RECT 186.480 14.865 186.760 15.145 ;
        RECT 188.265 14.865 188.545 15.145 ;
        RECT 191.120 14.865 191.400 15.145 ;
        RECT 192.905 14.865 193.185 15.145 ;
        RECT 177.200 14.205 177.480 14.485 ;
        RECT 178.985 14.205 179.265 14.485 ;
        RECT 181.840 14.205 182.120 14.485 ;
        RECT 183.625 14.205 183.905 14.485 ;
        RECT 186.480 14.205 186.760 14.485 ;
        RECT 188.265 14.205 188.545 14.485 ;
        RECT 191.120 14.205 191.400 14.485 ;
        RECT 192.905 14.205 193.185 14.485 ;
        RECT 177.200 13.545 177.480 13.825 ;
        RECT 178.985 13.545 179.265 13.825 ;
        RECT 181.840 13.545 182.120 13.825 ;
        RECT 183.625 13.545 183.905 13.825 ;
        RECT 186.480 13.545 186.760 13.825 ;
        RECT 188.265 13.545 188.545 13.825 ;
        RECT 191.120 13.545 191.400 13.825 ;
        RECT 192.905 13.545 193.185 13.825 ;
        RECT 177.200 12.885 177.480 13.165 ;
        RECT 178.985 12.885 179.265 13.165 ;
        RECT 181.840 12.885 182.120 13.165 ;
        RECT 183.625 12.885 183.905 13.165 ;
        RECT 186.480 12.885 186.760 13.165 ;
        RECT 188.265 12.885 188.545 13.165 ;
        RECT 191.120 12.885 191.400 13.165 ;
        RECT 192.905 12.885 193.185 13.165 ;
        RECT 177.200 12.225 177.480 12.505 ;
        RECT 178.985 12.225 179.265 12.505 ;
        RECT 181.840 12.225 182.120 12.505 ;
        RECT 183.625 12.225 183.905 12.505 ;
        RECT 186.480 12.225 186.760 12.505 ;
        RECT 188.265 12.225 188.545 12.505 ;
        RECT 191.120 12.225 191.400 12.505 ;
        RECT 192.905 12.225 193.185 12.505 ;
        RECT 177.200 11.565 177.480 11.845 ;
        RECT 178.985 11.565 179.265 11.845 ;
        RECT 181.840 11.565 182.120 11.845 ;
        RECT 183.625 11.565 183.905 11.845 ;
        RECT 186.480 11.565 186.760 11.845 ;
        RECT 188.265 11.565 188.545 11.845 ;
        RECT 191.120 11.565 191.400 11.845 ;
        RECT 192.905 11.565 193.185 11.845 ;
        RECT 177.200 10.905 177.480 11.185 ;
        RECT 178.985 10.905 179.265 11.185 ;
        RECT 181.840 10.905 182.120 11.185 ;
        RECT 183.625 10.905 183.905 11.185 ;
        RECT 186.480 10.905 186.760 11.185 ;
        RECT 188.265 10.905 188.545 11.185 ;
        RECT 191.120 10.905 191.400 11.185 ;
        RECT 192.905 10.905 193.185 11.185 ;
        RECT 177.200 10.245 177.480 10.525 ;
        RECT 178.985 10.245 179.265 10.525 ;
        RECT 181.840 10.245 182.120 10.525 ;
        RECT 183.625 10.245 183.905 10.525 ;
        RECT 186.480 10.245 186.760 10.525 ;
        RECT 188.265 10.245 188.545 10.525 ;
        RECT 191.120 10.245 191.400 10.525 ;
        RECT 192.905 10.245 193.185 10.525 ;
        RECT 177.200 9.585 177.480 9.865 ;
        RECT 178.985 9.585 179.265 9.865 ;
        RECT 181.840 9.585 182.120 9.865 ;
        RECT 183.625 9.585 183.905 9.865 ;
        RECT 186.480 9.585 186.760 9.865 ;
        RECT 188.265 9.585 188.545 9.865 ;
        RECT 191.120 9.585 191.400 9.865 ;
        RECT 192.905 9.585 193.185 9.865 ;
        RECT 177.200 8.925 177.480 9.205 ;
        RECT 178.985 8.925 179.265 9.205 ;
        RECT 181.840 8.925 182.120 9.205 ;
        RECT 183.625 8.925 183.905 9.205 ;
        RECT 186.480 8.925 186.760 9.205 ;
        RECT 188.265 8.925 188.545 9.205 ;
        RECT 191.120 8.925 191.400 9.205 ;
        RECT 192.905 8.925 193.185 9.205 ;
        RECT 4.660 8.140 4.940 8.420 ;
        RECT 22.850 8.140 23.130 8.420 ;
        RECT 42.160 8.140 42.440 8.420 ;
        RECT 56.990 8.140 57.270 8.420 ;
        RECT 4.660 7.480 4.940 7.760 ;
        RECT 22.850 7.480 23.130 7.760 ;
        RECT 42.160 7.480 42.440 7.760 ;
        RECT 56.990 7.480 57.270 7.760 ;
        RECT 4.660 6.820 4.940 7.100 ;
        RECT 22.850 6.820 23.130 7.100 ;
        RECT 42.160 6.820 42.440 7.100 ;
        RECT 56.990 6.820 57.270 7.100 ;
        RECT 0.900 4.740 1.180 5.020 ;
        RECT 2.040 4.740 2.320 5.020 ;
        RECT 8.080 4.770 8.360 5.050 ;
        RECT 8.740 4.770 9.020 5.050 ;
        RECT 9.400 4.770 9.680 5.050 ;
        RECT 14.610 4.740 14.890 5.020 ;
        RECT 15.270 4.740 15.550 5.020 ;
        RECT 15.930 4.740 16.210 5.020 ;
        RECT 17.970 4.740 18.250 5.020 ;
        RECT 18.630 4.740 18.910 5.020 ;
        RECT 19.290 4.740 19.570 5.020 ;
        RECT 26.270 4.770 26.550 5.050 ;
        RECT 26.930 4.770 27.210 5.050 ;
        RECT 27.590 4.770 27.870 5.050 ;
        RECT 32.800 4.740 33.080 5.020 ;
        RECT 33.460 4.740 33.740 5.020 ;
        RECT 34.120 4.740 34.400 5.020 ;
        RECT 36.160 4.740 36.440 5.020 ;
        RECT 36.820 4.740 37.100 5.020 ;
        RECT 37.480 4.740 37.760 5.020 ;
        RECT 39.540 4.740 39.820 5.020 ;
        RECT 45.580 4.770 45.860 5.050 ;
        RECT 46.240 4.770 46.520 5.050 ;
        RECT 46.900 4.770 47.180 5.050 ;
        RECT 52.110 4.740 52.390 5.020 ;
        RECT 52.770 4.740 53.050 5.020 ;
        RECT 53.430 4.740 53.710 5.020 ;
        RECT 60.410 4.770 60.690 5.050 ;
        RECT 61.070 4.770 61.350 5.050 ;
        RECT 61.730 4.770 62.010 5.050 ;
        RECT 66.940 4.740 67.220 5.020 ;
        RECT 67.600 4.740 67.880 5.020 ;
        RECT 68.260 4.740 68.540 5.020 ;
        RECT 70.300 4.740 70.580 5.020 ;
        RECT 70.960 4.740 71.240 5.020 ;
        RECT 71.620 4.740 71.900 5.020 ;
        RECT 73.680 4.740 73.960 5.020 ;
        RECT 74.680 4.740 74.960 5.020 ;
        RECT 75.340 4.740 75.620 5.020 ;
        RECT 76.000 4.740 76.280 5.020 ;
        RECT 76.920 4.740 77.200 5.020 ;
        RECT 77.580 4.740 77.860 5.020 ;
        RECT 78.240 4.740 78.520 5.020 ;
        RECT 79.260 4.740 79.540 5.020 ;
        RECT 79.920 4.740 80.200 5.020 ;
        RECT 80.580 4.740 80.860 5.020 ;
        RECT 82.520 4.740 82.800 5.020 ;
        RECT 83.180 4.740 83.460 5.020 ;
        RECT 83.840 4.740 84.120 5.020 ;
        RECT 84.760 4.740 85.040 5.020 ;
        RECT 85.420 4.740 85.700 5.020 ;
        RECT 86.080 4.740 86.360 5.020 ;
        RECT 87.000 4.740 87.280 5.020 ;
        RECT 87.660 4.740 87.940 5.020 ;
        RECT 88.320 4.740 88.600 5.020 ;
        RECT 89.240 4.740 89.520 5.020 ;
        RECT 89.900 4.740 90.180 5.020 ;
        RECT 90.560 4.740 90.840 5.020 ;
        RECT 91.480 4.740 91.760 5.020 ;
        RECT 92.140 4.740 92.420 5.020 ;
        RECT 92.800 4.740 93.080 5.020 ;
        RECT 93.840 4.740 94.120 5.020 ;
        RECT 94.840 4.740 95.120 5.020 ;
        RECT 95.500 4.740 95.780 5.020 ;
        RECT 96.160 4.740 96.440 5.020 ;
        RECT 97.080 4.740 97.360 5.020 ;
        RECT 97.740 4.740 98.020 5.020 ;
        RECT 98.400 4.740 98.680 5.020 ;
        RECT 99.320 4.740 99.600 5.020 ;
        RECT 99.980 4.740 100.260 5.020 ;
        RECT 100.640 4.740 100.920 5.020 ;
        RECT 101.660 4.740 101.940 5.020 ;
        RECT 102.320 4.740 102.600 5.020 ;
        RECT 102.980 4.740 103.260 5.020 ;
        RECT 104.920 4.740 105.200 5.020 ;
        RECT 105.580 4.740 105.860 5.020 ;
        RECT 106.240 4.740 106.520 5.020 ;
        RECT 107.160 4.740 107.440 5.020 ;
        RECT 107.820 4.740 108.100 5.020 ;
        RECT 108.480 4.740 108.760 5.020 ;
        RECT 109.400 4.740 109.680 5.020 ;
        RECT 110.060 4.740 110.340 5.020 ;
        RECT 110.720 4.740 111.000 5.020 ;
        RECT 111.640 4.740 111.920 5.020 ;
        RECT 112.300 4.740 112.580 5.020 ;
        RECT 112.960 4.740 113.240 5.020 ;
        RECT 114.000 4.740 114.280 5.020 ;
        RECT 115.000 4.740 115.280 5.020 ;
        RECT 115.660 4.740 115.940 5.020 ;
        RECT 116.320 4.740 116.600 5.020 ;
        RECT 117.240 4.740 117.520 5.020 ;
        RECT 117.900 4.740 118.180 5.020 ;
        RECT 118.560 4.740 118.840 5.020 ;
        RECT 119.480 4.740 119.760 5.020 ;
        RECT 120.140 4.740 120.420 5.020 ;
        RECT 120.800 4.740 121.080 5.020 ;
        RECT 121.820 4.740 122.100 5.020 ;
        RECT 122.480 4.740 122.760 5.020 ;
        RECT 123.140 4.740 123.420 5.020 ;
        RECT 125.080 4.740 125.360 5.020 ;
        RECT 125.740 4.740 126.020 5.020 ;
        RECT 126.400 4.740 126.680 5.020 ;
        RECT 127.320 4.740 127.600 5.020 ;
        RECT 127.980 4.740 128.260 5.020 ;
        RECT 128.640 4.740 128.920 5.020 ;
        RECT 129.560 4.740 129.840 5.020 ;
        RECT 130.220 4.740 130.500 5.020 ;
        RECT 130.880 4.740 131.160 5.020 ;
        RECT 131.800 4.740 132.080 5.020 ;
        RECT 132.460 4.740 132.740 5.020 ;
        RECT 133.120 4.740 133.400 5.020 ;
        RECT 134.160 4.740 134.440 5.020 ;
        RECT 135.160 4.740 135.440 5.020 ;
        RECT 135.820 4.740 136.100 5.020 ;
        RECT 136.480 4.740 136.760 5.020 ;
        RECT 137.400 4.740 137.680 5.020 ;
        RECT 138.060 4.740 138.340 5.020 ;
        RECT 138.720 4.740 139.000 5.020 ;
        RECT 139.640 4.740 139.920 5.020 ;
        RECT 140.300 4.740 140.580 5.020 ;
        RECT 140.960 4.740 141.240 5.020 ;
        RECT 141.880 4.740 142.160 5.020 ;
        RECT 142.540 4.740 142.820 5.020 ;
        RECT 143.200 4.740 143.480 5.020 ;
        RECT 144.220 4.740 144.500 5.020 ;
        RECT 144.880 4.740 145.160 5.020 ;
        RECT 145.540 4.740 145.820 5.020 ;
        RECT 147.480 4.740 147.760 5.020 ;
        RECT 148.140 4.740 148.420 5.020 ;
        RECT 148.800 4.740 149.080 5.020 ;
        RECT 149.720 4.740 150.000 5.020 ;
        RECT 150.380 4.740 150.660 5.020 ;
        RECT 151.040 4.740 151.320 5.020 ;
        RECT 151.960 4.740 152.240 5.020 ;
        RECT 152.620 4.740 152.900 5.020 ;
        RECT 153.280 4.740 153.560 5.020 ;
        RECT 154.320 4.740 154.600 5.020 ;
        RECT 155.320 4.740 155.600 5.020 ;
        RECT 155.980 4.740 156.260 5.020 ;
        RECT 156.640 4.740 156.920 5.020 ;
        RECT 157.560 4.740 157.840 5.020 ;
        RECT 158.220 4.740 158.500 5.020 ;
        RECT 158.880 4.740 159.160 5.020 ;
        RECT 159.800 4.740 160.080 5.020 ;
        RECT 160.460 4.740 160.740 5.020 ;
        RECT 161.120 4.740 161.400 5.020 ;
        RECT 162.040 4.740 162.320 5.020 ;
        RECT 162.700 4.740 162.980 5.020 ;
        RECT 163.360 4.740 163.640 5.020 ;
        RECT 164.280 4.740 164.560 5.020 ;
        RECT 164.940 4.740 165.220 5.020 ;
        RECT 165.600 4.740 165.880 5.020 ;
        RECT 166.620 4.740 166.900 5.020 ;
        RECT 167.280 4.740 167.560 5.020 ;
        RECT 167.940 4.740 168.220 5.020 ;
        RECT 169.880 4.740 170.160 5.020 ;
        RECT 170.540 4.740 170.820 5.020 ;
        RECT 171.200 4.740 171.480 5.020 ;
        RECT 172.120 4.740 172.400 5.020 ;
        RECT 172.780 4.740 173.060 5.020 ;
        RECT 173.440 4.740 173.720 5.020 ;
        RECT 174.460 4.740 174.740 5.020 ;
        RECT 0.900 0.820 1.180 1.100 ;
        RECT 2.040 0.820 2.320 1.100 ;
        RECT 7.480 0.820 7.760 1.100 ;
        RECT 8.140 0.820 8.420 1.100 ;
        RECT 8.800 0.820 9.080 1.100 ;
        RECT 14.350 0.820 14.630 1.100 ;
        RECT 15.670 0.820 15.950 1.100 ;
        RECT 17.710 0.820 17.990 1.100 ;
        RECT 19.030 0.820 19.310 1.100 ;
        RECT 25.670 0.820 25.950 1.100 ;
        RECT 26.330 0.820 26.610 1.100 ;
        RECT 26.990 0.820 27.270 1.100 ;
        RECT 32.540 0.820 32.820 1.100 ;
        RECT 33.860 0.820 34.140 1.100 ;
        RECT 35.900 0.820 36.180 1.100 ;
        RECT 37.220 0.820 37.500 1.100 ;
        RECT 39.540 0.820 39.820 1.100 ;
        RECT 44.980 0.820 45.260 1.100 ;
        RECT 45.640 0.820 45.920 1.100 ;
        RECT 46.300 0.820 46.580 1.100 ;
        RECT 51.850 0.820 52.130 1.100 ;
        RECT 53.170 0.820 53.450 1.100 ;
        RECT 59.810 0.820 60.090 1.100 ;
        RECT 60.470 0.820 60.750 1.100 ;
        RECT 61.130 0.820 61.410 1.100 ;
        RECT 66.680 0.820 66.960 1.100 ;
        RECT 68.000 0.820 68.280 1.100 ;
        RECT 70.040 0.820 70.320 1.100 ;
        RECT 71.360 0.820 71.640 1.100 ;
        RECT 73.680 0.820 73.960 1.100 ;
        RECT 74.680 0.820 74.960 1.100 ;
        RECT 75.340 0.820 75.620 1.100 ;
        RECT 76.000 0.820 76.280 1.100 ;
        RECT 76.920 0.820 77.200 1.100 ;
        RECT 77.580 0.820 77.860 1.100 ;
        RECT 78.240 0.820 78.520 1.100 ;
        RECT 79.000 0.820 79.280 1.100 ;
        RECT 80.320 0.820 80.600 1.100 ;
        RECT 82.520 0.820 82.800 1.100 ;
        RECT 83.180 0.820 83.460 1.100 ;
        RECT 83.840 0.820 84.120 1.100 ;
        RECT 84.760 0.820 85.040 1.100 ;
        RECT 85.420 0.820 85.700 1.100 ;
        RECT 86.080 0.820 86.360 1.100 ;
        RECT 87.000 0.820 87.280 1.100 ;
        RECT 87.660 0.820 87.940 1.100 ;
        RECT 88.320 0.820 88.600 1.100 ;
        RECT 89.240 0.820 89.520 1.100 ;
        RECT 89.900 0.820 90.180 1.100 ;
        RECT 90.560 0.820 90.840 1.100 ;
        RECT 91.480 0.820 91.760 1.100 ;
        RECT 92.140 0.820 92.420 1.100 ;
        RECT 92.800 0.820 93.080 1.100 ;
        RECT 93.840 0.820 94.120 1.100 ;
        RECT 94.840 0.820 95.120 1.100 ;
        RECT 95.500 0.820 95.780 1.100 ;
        RECT 96.160 0.820 96.440 1.100 ;
        RECT 97.080 0.820 97.360 1.100 ;
        RECT 97.740 0.820 98.020 1.100 ;
        RECT 98.400 0.820 98.680 1.100 ;
        RECT 99.320 0.820 99.600 1.100 ;
        RECT 99.980 0.820 100.260 1.100 ;
        RECT 100.640 0.820 100.920 1.100 ;
        RECT 101.400 0.820 101.680 1.100 ;
        RECT 102.720 0.820 103.000 1.100 ;
        RECT 104.920 0.820 105.200 1.100 ;
        RECT 105.580 0.820 105.860 1.100 ;
        RECT 106.240 0.820 106.520 1.100 ;
        RECT 107.160 0.820 107.440 1.100 ;
        RECT 107.820 0.820 108.100 1.100 ;
        RECT 108.480 0.820 108.760 1.100 ;
        RECT 109.400 0.820 109.680 1.100 ;
        RECT 110.060 0.820 110.340 1.100 ;
        RECT 110.720 0.820 111.000 1.100 ;
        RECT 111.640 0.820 111.920 1.100 ;
        RECT 112.300 0.820 112.580 1.100 ;
        RECT 112.960 0.820 113.240 1.100 ;
        RECT 114.000 0.820 114.280 1.100 ;
        RECT 115.000 0.820 115.280 1.100 ;
        RECT 115.660 0.820 115.940 1.100 ;
        RECT 116.320 0.820 116.600 1.100 ;
        RECT 117.240 0.820 117.520 1.100 ;
        RECT 117.900 0.820 118.180 1.100 ;
        RECT 118.560 0.820 118.840 1.100 ;
        RECT 119.480 0.820 119.760 1.100 ;
        RECT 120.140 0.820 120.420 1.100 ;
        RECT 120.800 0.820 121.080 1.100 ;
        RECT 121.560 0.820 121.840 1.100 ;
        RECT 122.880 0.820 123.160 1.100 ;
        RECT 125.080 0.820 125.360 1.100 ;
        RECT 125.740 0.820 126.020 1.100 ;
        RECT 126.400 0.820 126.680 1.100 ;
        RECT 127.320 0.820 127.600 1.100 ;
        RECT 127.980 0.820 128.260 1.100 ;
        RECT 128.640 0.820 128.920 1.100 ;
        RECT 129.560 0.820 129.840 1.100 ;
        RECT 130.220 0.820 130.500 1.100 ;
        RECT 130.880 0.820 131.160 1.100 ;
        RECT 131.800 0.820 132.080 1.100 ;
        RECT 132.460 0.820 132.740 1.100 ;
        RECT 133.120 0.820 133.400 1.100 ;
        RECT 134.160 0.820 134.440 1.100 ;
        RECT 135.160 0.820 135.440 1.100 ;
        RECT 135.820 0.820 136.100 1.100 ;
        RECT 136.480 0.820 136.760 1.100 ;
        RECT 137.400 0.820 137.680 1.100 ;
        RECT 138.060 0.820 138.340 1.100 ;
        RECT 138.720 0.820 139.000 1.100 ;
        RECT 139.640 0.820 139.920 1.100 ;
        RECT 140.300 0.820 140.580 1.100 ;
        RECT 140.960 0.820 141.240 1.100 ;
        RECT 141.880 0.820 142.160 1.100 ;
        RECT 142.540 0.820 142.820 1.100 ;
        RECT 143.200 0.820 143.480 1.100 ;
        RECT 143.960 0.820 144.240 1.100 ;
        RECT 145.280 0.820 145.560 1.100 ;
        RECT 147.480 0.820 147.760 1.100 ;
        RECT 148.140 0.820 148.420 1.100 ;
        RECT 148.800 0.820 149.080 1.100 ;
        RECT 149.720 0.820 150.000 1.100 ;
        RECT 150.380 0.820 150.660 1.100 ;
        RECT 151.040 0.820 151.320 1.100 ;
        RECT 151.960 0.820 152.240 1.100 ;
        RECT 152.620 0.820 152.900 1.100 ;
        RECT 153.280 0.820 153.560 1.100 ;
        RECT 154.320 0.820 154.600 1.100 ;
        RECT 155.320 0.820 155.600 1.100 ;
        RECT 155.980 0.820 156.260 1.100 ;
        RECT 156.640 0.820 156.920 1.100 ;
        RECT 157.560 0.820 157.840 1.100 ;
        RECT 158.220 0.820 158.500 1.100 ;
        RECT 158.880 0.820 159.160 1.100 ;
        RECT 159.800 0.820 160.080 1.100 ;
        RECT 160.460 0.820 160.740 1.100 ;
        RECT 161.120 0.820 161.400 1.100 ;
        RECT 162.040 0.820 162.320 1.100 ;
        RECT 162.700 0.820 162.980 1.100 ;
        RECT 163.360 0.820 163.640 1.100 ;
        RECT 164.280 0.820 164.560 1.100 ;
        RECT 164.940 0.820 165.220 1.100 ;
        RECT 165.600 0.820 165.880 1.100 ;
        RECT 166.360 0.820 166.640 1.100 ;
        RECT 167.680 0.820 167.960 1.100 ;
        RECT 169.880 0.820 170.160 1.100 ;
        RECT 170.540 0.820 170.820 1.100 ;
        RECT 171.200 0.820 171.480 1.100 ;
        RECT 172.120 0.820 172.400 1.100 ;
        RECT 172.780 0.820 173.060 1.100 ;
        RECT 173.440 0.820 173.720 1.100 ;
        RECT 174.460 0.820 174.740 1.100 ;
      LAYER Metal4 ;
        RECT 4.610 47.805 4.990 48.185 ;
        RECT 4.635 47.525 4.965 47.805 ;
        RECT 4.610 47.145 4.990 47.525 ;
        RECT 4.635 46.865 4.965 47.145 ;
        RECT 4.610 46.485 4.990 46.865 ;
        RECT 4.635 8.470 4.965 46.485 ;
        RECT 56.940 45.105 57.320 45.485 ;
        RECT 56.965 44.825 57.295 45.105 ;
        RECT 56.940 44.445 57.320 44.825 ;
        RECT 56.965 44.165 57.295 44.445 ;
        RECT 56.940 43.785 57.320 44.165 ;
        RECT 42.110 24.905 42.490 25.285 ;
        RECT 42.135 24.625 42.465 24.905 ;
        RECT 42.110 24.245 42.490 24.625 ;
        RECT 42.135 23.965 42.465 24.245 ;
        RECT 42.110 23.585 42.490 23.965 ;
        RECT 22.800 22.205 23.180 22.585 ;
        RECT 22.825 21.925 23.155 22.205 ;
        RECT 22.800 21.545 23.180 21.925 ;
        RECT 22.825 21.265 23.155 21.545 ;
        RECT 22.800 20.885 23.180 21.265 ;
        RECT 22.825 8.470 23.155 20.885 ;
        RECT 42.135 8.470 42.465 23.585 ;
        RECT 56.965 8.470 57.295 43.785 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 42.110 8.090 42.490 8.470 ;
        RECT 56.940 8.090 57.320 8.470 ;
        RECT 4.635 7.810 4.965 8.090 ;
        RECT 22.825 7.810 23.155 8.090 ;
        RECT 42.135 7.810 42.465 8.090 ;
        RECT 56.965 7.810 57.295 8.090 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 42.110 7.430 42.490 7.810 ;
        RECT 56.940 7.430 57.320 7.810 ;
        RECT 4.635 7.150 4.965 7.430 ;
        RECT 22.825 7.150 23.155 7.430 ;
        RECT 42.135 7.150 42.465 7.430 ;
        RECT 56.965 7.150 57.295 7.430 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 42.110 6.770 42.490 7.150 ;
        RECT 56.940 6.770 57.320 7.150 ;
  END
END efuse_array
END LIBRARY

