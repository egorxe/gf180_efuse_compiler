module efuse_array(nPRESET, SENSE, COL_PROG, LINE, DO);
  output [7:0] DO;
  wire [7:0] DO;
  input [7:0] COL_PROG;
  wire [7:0] COL_PROG;
  input [15:0] LINE;
  wire [15:0] LINE;
  input SENSE;
  wire SENSE;
  input nPRESET;
  wire nPRESET;
endmodule

