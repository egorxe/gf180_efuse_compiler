VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array
  CLASS BLOCK ;
  FOREIGN efuse_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 717.540 BY 60.305 ;
  PIN COL_PROG[0]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 683.600 59.415 683.940 60.305 ;
    END
  END COL_PROG[0]
  PIN COL_PROG[1]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 688.240 59.415 688.580 60.305 ;
    END
  END COL_PROG[1]
  PIN COL_PROG[2]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 692.880 59.415 693.220 60.305 ;
    END
  END COL_PROG[2]
  PIN COL_PROG[3]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 697.520 59.415 697.860 60.305 ;
    END
  END COL_PROG[3]
  PIN COL_PROG[4]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 702.160 59.415 702.500 60.305 ;
    END
  END COL_PROG[4]
  PIN COL_PROG[5]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 706.800 59.415 707.140 60.305 ;
    END
  END COL_PROG[5]
  PIN COL_PROG[6]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 711.440 59.415 711.780 60.305 ;
    END
  END COL_PROG[6]
  PIN COL_PROG[7]
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER Metal1 ;
        RECT 716.080 59.415 716.420 60.305 ;
    END
  END COL_PROG[7]
  PIN DO[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.720 1.770 17.100 2.150 ;
        RECT 16.745 0.000 17.075 1.770 ;
    END
  END DO[0]
  PIN LINE[0]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 18.305 2.770 18.685 3.150 ;
        RECT 18.330 0.000 18.660 2.770 ;
    END
  END LINE[0]
  PIN DO[1]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.910 1.770 35.290 2.150 ;
        RECT 34.935 0.000 35.265 1.770 ;
    END
  END DO[1]
  PIN DO[2]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.860 1.770 51.240 2.150 ;
        RECT 50.885 0.000 51.215 1.770 ;
    END
  END DO[2]
  PIN DO[3]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 65.690 1.770 66.070 2.150 ;
        RECT 65.715 0.000 66.045 1.770 ;
    END
  END DO[3]
  PIN LINE[1]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 67.275 2.770 67.655 3.150 ;
        RECT 67.300 0.000 67.630 2.770 ;
    END
  END LINE[1]
  PIN DO[4]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.000 1.770 85.380 2.150 ;
        RECT 85.025 0.000 85.355 1.770 ;
    END
  END DO[4]
  PIN DO[5]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 99.830 1.770 100.210 2.150 ;
        RECT 99.855 0.000 100.185 1.770 ;
    END
  END DO[5]
  PIN LINE[2]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 101.415 2.770 101.795 3.150 ;
        RECT 101.440 0.000 101.770 2.770 ;
    END
  END LINE[2]
  PIN DO[6]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 119.140 1.770 119.520 2.150 ;
        RECT 119.165 0.000 119.495 1.770 ;
    END
  END DO[6]
  PIN DO[7]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.970 1.770 134.350 2.150 ;
        RECT 133.995 0.000 134.325 1.770 ;
    END
  END DO[7]
  PIN LINE[3]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 141.155 2.770 141.535 3.150 ;
        RECT 141.180 0.000 141.510 2.770 ;
    END
  END LINE[3]
  PIN LINE[4]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 182.595 2.770 182.975 3.150 ;
        RECT 182.620 0.000 182.950 2.770 ;
    END
  END LINE[4]
  PIN LINE[5]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 226.275 2.770 226.655 3.150 ;
        RECT 226.300 0.000 226.630 2.770 ;
    END
  END LINE[5]
  PIN LINE[6]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 267.715 2.770 268.095 3.150 ;
        RECT 267.740 0.000 268.070 2.770 ;
    END
  END LINE[6]
  PIN LINE[7]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 311.395 2.770 311.775 3.150 ;
        RECT 311.420 0.000 311.750 2.770 ;
    END
  END LINE[7]
  PIN LINE[8]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 352.835 2.770 353.215 3.150 ;
        RECT 352.860 0.000 353.190 2.770 ;
    END
  END LINE[8]
  PIN LINE[9]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 396.515 2.770 396.895 3.150 ;
        RECT 396.540 0.000 396.870 2.770 ;
    END
  END LINE[9]
  PIN LINE[10]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 437.955 2.770 438.335 3.150 ;
        RECT 437.980 0.000 438.310 2.770 ;
    END
  END LINE[10]
  PIN LINE[11]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 481.635 2.770 482.015 3.150 ;
        RECT 481.660 0.000 481.990 2.770 ;
    END
  END LINE[11]
  PIN LINE[12]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 523.075 2.770 523.455 3.150 ;
        RECT 523.100 0.000 523.430 2.770 ;
    END
  END LINE[12]
  PIN LINE[13]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 566.755 2.770 567.135 3.150 ;
        RECT 566.780 0.000 567.110 2.770 ;
    END
  END LINE[13]
  PIN LINE[14]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 608.195 2.770 608.575 3.150 ;
        RECT 608.220 0.000 608.550 2.770 ;
    END
  END LINE[14]
  PIN LINE[15]
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal2 ;
        RECT 651.875 2.770 652.255 3.150 ;
        RECT 651.900 0.000 652.230 2.770 ;
    END
  END LINE[15]
  PIN SENSE
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER Metal3 ;
        RECT 4.170 3.775 4.550 3.800 ;
        RECT 22.360 3.775 22.740 3.800 ;
        RECT 38.310 3.775 38.690 3.800 ;
        RECT 53.140 3.775 53.520 3.800 ;
        RECT 72.450 3.775 72.830 3.800 ;
        RECT 87.280 3.775 87.660 3.800 ;
        RECT 106.590 3.775 106.970 3.800 ;
        RECT 121.420 3.775 121.800 3.800 ;
        RECT 4.170 3.445 121.800 3.775 ;
        RECT 4.170 3.420 4.550 3.445 ;
        RECT 22.360 3.420 22.740 3.445 ;
        RECT 38.310 3.420 38.690 3.445 ;
        RECT 53.140 3.420 53.520 3.445 ;
        RECT 72.450 3.420 72.830 3.445 ;
        RECT 87.280 3.420 87.660 3.445 ;
        RECT 106.590 3.420 106.970 3.445 ;
        RECT 121.420 3.420 121.800 3.445 ;
    END
  END SENSE
  PIN nPRESET
    ANTENNAGATEAREA 7.600000 ;
    PORT
      LAYER Metal3 ;
        RECT 4.580 3.115 4.960 3.140 ;
        RECT 22.770 3.115 23.150 3.140 ;
        RECT 38.720 3.115 39.100 3.140 ;
        RECT 53.550 3.115 53.930 3.140 ;
        RECT 72.860 3.115 73.240 3.140 ;
        RECT 87.690 3.115 88.070 3.140 ;
        RECT 107.000 3.115 107.380 3.140 ;
        RECT 121.830 3.115 122.210 3.140 ;
        RECT 4.580 2.785 122.210 3.115 ;
        RECT 4.580 2.760 4.960 2.785 ;
        RECT 22.770 2.760 23.150 2.785 ;
        RECT 38.720 2.760 39.100 2.785 ;
        RECT 53.550 2.760 53.930 2.785 ;
        RECT 72.860 2.760 73.240 2.785 ;
        RECT 87.690 2.760 88.070 2.785 ;
        RECT 107.000 2.760 107.380 2.785 ;
        RECT 121.830 2.760 122.210 2.785 ;
    END
  END nPRESET
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 0.000 57.805 717.540 60.305 ;
        RECT 0.000 49.035 1.910 57.805 ;
        RECT 10.290 49.035 12.200 57.805 ;
        RECT 20.575 49.035 22.485 57.805 ;
        RECT 30.865 49.035 32.775 57.805 ;
        RECT 41.150 49.035 44.480 57.805 ;
        RECT 52.860 49.035 54.770 57.805 ;
        RECT 63.145 49.035 65.055 57.805 ;
        RECT 73.435 49.035 75.345 57.805 ;
        RECT 83.720 49.035 87.050 57.805 ;
        RECT 95.430 49.035 97.340 57.805 ;
        RECT 105.715 49.035 107.625 57.805 ;
        RECT 116.005 49.035 117.915 57.805 ;
        RECT 126.290 49.035 129.620 57.805 ;
        RECT 138.000 49.035 139.910 57.805 ;
        RECT 148.285 49.035 150.195 57.805 ;
        RECT 158.575 49.035 160.485 57.805 ;
        RECT 168.860 49.035 172.190 57.805 ;
        RECT 180.570 49.035 182.480 57.805 ;
        RECT 190.855 49.035 192.765 57.805 ;
        RECT 201.145 49.035 203.055 57.805 ;
        RECT 211.430 49.035 214.760 57.805 ;
        RECT 223.140 49.035 225.050 57.805 ;
        RECT 233.425 49.035 235.335 57.805 ;
        RECT 243.715 49.035 245.625 57.805 ;
        RECT 254.000 49.035 257.330 57.805 ;
        RECT 265.710 49.035 267.620 57.805 ;
        RECT 275.995 49.035 277.905 57.805 ;
        RECT 286.285 49.035 288.195 57.805 ;
        RECT 296.570 49.035 299.900 57.805 ;
        RECT 308.280 49.035 310.190 57.805 ;
        RECT 318.565 49.035 320.475 57.805 ;
        RECT 328.855 49.035 330.765 57.805 ;
        RECT 339.140 49.035 342.470 57.805 ;
        RECT 350.850 49.035 352.760 57.805 ;
        RECT 361.135 49.035 363.045 57.805 ;
        RECT 371.425 49.035 373.335 57.805 ;
        RECT 381.710 49.035 385.040 57.805 ;
        RECT 393.420 49.035 395.330 57.805 ;
        RECT 403.705 49.035 405.615 57.805 ;
        RECT 413.995 49.035 415.905 57.805 ;
        RECT 424.280 49.035 427.610 57.805 ;
        RECT 435.990 49.035 437.900 57.805 ;
        RECT 446.275 49.035 448.185 57.805 ;
        RECT 456.565 49.035 458.475 57.805 ;
        RECT 466.850 49.035 470.180 57.805 ;
        RECT 478.560 49.035 480.470 57.805 ;
        RECT 488.845 49.035 490.755 57.805 ;
        RECT 499.135 49.035 501.045 57.805 ;
        RECT 509.420 49.035 512.750 57.805 ;
        RECT 521.130 49.035 523.040 57.805 ;
        RECT 531.415 49.035 533.325 57.805 ;
        RECT 541.705 49.035 543.615 57.805 ;
        RECT 551.990 49.035 555.320 57.805 ;
        RECT 563.700 49.035 565.610 57.805 ;
        RECT 573.985 49.035 575.895 57.805 ;
        RECT 584.275 49.035 586.185 57.805 ;
        RECT 594.560 49.035 597.890 57.805 ;
        RECT 606.270 49.035 608.180 57.805 ;
        RECT 616.555 49.035 618.465 57.805 ;
        RECT 626.845 49.035 628.755 57.805 ;
        RECT 637.130 49.035 640.460 57.805 ;
        RECT 648.840 49.035 650.750 57.805 ;
        RECT 659.125 49.035 661.035 57.805 ;
        RECT 669.415 49.035 671.325 57.805 ;
        RECT 678.620 49.035 681.610 57.805 ;
        RECT 678.620 6.470 681.120 49.035 ;
        RECT 0.000 3.970 681.120 6.470 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 682.335 55.495 684.450 55.805 ;
        RECT 686.975 55.495 689.090 55.805 ;
        RECT 691.615 55.495 693.730 55.805 ;
        RECT 696.255 55.495 698.370 55.805 ;
        RECT 700.895 55.495 703.010 55.805 ;
        RECT 705.535 55.495 707.650 55.805 ;
        RECT 710.175 55.495 712.290 55.805 ;
        RECT 714.815 55.495 716.930 55.805 ;
        RECT 682.310 55.115 684.475 55.495 ;
        RECT 686.950 55.115 689.115 55.495 ;
        RECT 691.590 55.115 693.755 55.495 ;
        RECT 696.230 55.115 698.395 55.495 ;
        RECT 700.870 55.115 703.035 55.495 ;
        RECT 705.510 55.115 707.675 55.495 ;
        RECT 710.150 55.115 712.315 55.495 ;
        RECT 714.790 55.115 716.955 55.495 ;
        RECT 682.335 54.835 684.450 55.115 ;
        RECT 686.975 54.835 689.090 55.115 ;
        RECT 691.615 54.835 693.730 55.115 ;
        RECT 696.255 54.835 698.370 55.115 ;
        RECT 700.895 54.835 703.010 55.115 ;
        RECT 705.535 54.835 707.650 55.115 ;
        RECT 710.175 54.835 712.290 55.115 ;
        RECT 714.815 54.835 716.930 55.115 ;
        RECT 682.310 54.455 684.475 54.835 ;
        RECT 686.950 54.455 689.115 54.835 ;
        RECT 691.590 54.455 693.755 54.835 ;
        RECT 696.230 54.455 698.395 54.835 ;
        RECT 700.870 54.455 703.035 54.835 ;
        RECT 705.510 54.455 707.675 54.835 ;
        RECT 710.150 54.455 712.315 54.835 ;
        RECT 714.790 54.455 716.955 54.835 ;
        RECT 682.335 54.175 684.450 54.455 ;
        RECT 686.975 54.175 689.090 54.455 ;
        RECT 691.615 54.175 693.730 54.455 ;
        RECT 696.255 54.175 698.370 54.455 ;
        RECT 700.895 54.175 703.010 54.455 ;
        RECT 705.535 54.175 707.650 54.455 ;
        RECT 710.175 54.175 712.290 54.455 ;
        RECT 714.815 54.175 716.930 54.455 ;
        RECT 682.310 53.795 684.475 54.175 ;
        RECT 686.950 53.795 689.115 54.175 ;
        RECT 691.590 53.795 693.755 54.175 ;
        RECT 696.230 53.795 698.395 54.175 ;
        RECT 700.870 53.795 703.035 54.175 ;
        RECT 705.510 53.795 707.675 54.175 ;
        RECT 710.150 53.795 712.315 54.175 ;
        RECT 714.790 53.795 716.955 54.175 ;
        RECT 682.335 53.515 684.450 53.795 ;
        RECT 686.975 53.515 689.090 53.795 ;
        RECT 691.615 53.515 693.730 53.795 ;
        RECT 696.255 53.515 698.370 53.795 ;
        RECT 700.895 53.515 703.010 53.795 ;
        RECT 705.535 53.515 707.650 53.795 ;
        RECT 710.175 53.515 712.290 53.795 ;
        RECT 714.815 53.515 716.930 53.795 ;
        RECT 682.310 53.135 684.475 53.515 ;
        RECT 686.950 53.135 689.115 53.515 ;
        RECT 691.590 53.135 693.755 53.515 ;
        RECT 696.230 53.135 698.395 53.515 ;
        RECT 700.870 53.135 703.035 53.515 ;
        RECT 705.510 53.135 707.675 53.515 ;
        RECT 710.150 53.135 712.315 53.515 ;
        RECT 714.790 53.135 716.955 53.515 ;
        RECT 682.335 52.855 684.450 53.135 ;
        RECT 686.975 52.855 689.090 53.135 ;
        RECT 691.615 52.855 693.730 53.135 ;
        RECT 696.255 52.855 698.370 53.135 ;
        RECT 700.895 52.855 703.010 53.135 ;
        RECT 705.535 52.855 707.650 53.135 ;
        RECT 710.175 52.855 712.290 53.135 ;
        RECT 714.815 52.855 716.930 53.135 ;
        RECT 682.310 52.475 684.475 52.855 ;
        RECT 686.950 52.475 689.115 52.855 ;
        RECT 691.590 52.475 693.755 52.855 ;
        RECT 696.230 52.475 698.395 52.855 ;
        RECT 700.870 52.475 703.035 52.855 ;
        RECT 705.510 52.475 707.675 52.855 ;
        RECT 710.150 52.475 712.315 52.855 ;
        RECT 714.790 52.475 716.955 52.855 ;
        RECT 682.335 52.195 684.450 52.475 ;
        RECT 686.975 52.195 689.090 52.475 ;
        RECT 691.615 52.195 693.730 52.475 ;
        RECT 696.255 52.195 698.370 52.475 ;
        RECT 700.895 52.195 703.010 52.475 ;
        RECT 705.535 52.195 707.650 52.475 ;
        RECT 710.175 52.195 712.290 52.475 ;
        RECT 714.815 52.195 716.930 52.475 ;
        RECT 682.310 51.815 684.475 52.195 ;
        RECT 686.950 51.815 689.115 52.195 ;
        RECT 691.590 51.815 693.755 52.195 ;
        RECT 696.230 51.815 698.395 52.195 ;
        RECT 700.870 51.815 703.035 52.195 ;
        RECT 705.510 51.815 707.675 52.195 ;
        RECT 710.150 51.815 712.315 52.195 ;
        RECT 714.790 51.815 716.955 52.195 ;
        RECT 682.335 51.535 684.450 51.815 ;
        RECT 686.975 51.535 689.090 51.815 ;
        RECT 691.615 51.535 693.730 51.815 ;
        RECT 696.255 51.535 698.370 51.815 ;
        RECT 700.895 51.535 703.010 51.815 ;
        RECT 705.535 51.535 707.650 51.815 ;
        RECT 710.175 51.535 712.290 51.815 ;
        RECT 714.815 51.535 716.930 51.815 ;
        RECT 682.310 51.155 684.475 51.535 ;
        RECT 686.950 51.155 689.115 51.535 ;
        RECT 691.590 51.155 693.755 51.535 ;
        RECT 696.230 51.155 698.395 51.535 ;
        RECT 700.870 51.155 703.035 51.535 ;
        RECT 705.510 51.155 707.675 51.535 ;
        RECT 710.150 51.155 712.315 51.535 ;
        RECT 714.790 51.155 716.955 51.535 ;
        RECT 682.335 50.875 684.450 51.155 ;
        RECT 686.975 50.875 689.090 51.155 ;
        RECT 691.615 50.875 693.730 51.155 ;
        RECT 696.255 50.875 698.370 51.155 ;
        RECT 700.895 50.875 703.010 51.155 ;
        RECT 705.535 50.875 707.650 51.155 ;
        RECT 710.175 50.875 712.290 51.155 ;
        RECT 714.815 50.875 716.930 51.155 ;
        RECT 682.310 50.495 684.475 50.875 ;
        RECT 686.950 50.495 689.115 50.875 ;
        RECT 691.590 50.495 693.755 50.875 ;
        RECT 696.230 50.495 698.395 50.875 ;
        RECT 700.870 50.495 703.035 50.875 ;
        RECT 705.510 50.495 707.675 50.875 ;
        RECT 710.150 50.495 712.315 50.875 ;
        RECT 714.790 50.495 716.955 50.875 ;
        RECT 682.335 18.495 684.450 50.495 ;
        RECT 686.975 18.495 689.090 50.495 ;
        RECT 691.615 18.495 693.730 50.495 ;
        RECT 696.255 18.495 698.370 50.495 ;
        RECT 700.895 18.495 703.010 50.495 ;
        RECT 705.535 18.495 707.650 50.495 ;
        RECT 710.175 18.495 712.290 50.495 ;
        RECT 714.815 18.495 716.930 50.495 ;
        RECT 682.310 18.115 684.475 18.495 ;
        RECT 686.950 18.115 689.115 18.495 ;
        RECT 691.590 18.115 693.755 18.495 ;
        RECT 696.230 18.115 698.395 18.495 ;
        RECT 700.870 18.115 703.035 18.495 ;
        RECT 705.510 18.115 707.675 18.495 ;
        RECT 710.150 18.115 712.315 18.495 ;
        RECT 714.790 18.115 716.955 18.495 ;
        RECT 682.335 17.835 684.450 18.115 ;
        RECT 686.975 17.835 689.090 18.115 ;
        RECT 691.615 17.835 693.730 18.115 ;
        RECT 696.255 17.835 698.370 18.115 ;
        RECT 700.895 17.835 703.010 18.115 ;
        RECT 705.535 17.835 707.650 18.115 ;
        RECT 710.175 17.835 712.290 18.115 ;
        RECT 714.815 17.835 716.930 18.115 ;
        RECT 682.310 17.455 684.475 17.835 ;
        RECT 686.950 17.455 689.115 17.835 ;
        RECT 691.590 17.455 693.755 17.835 ;
        RECT 696.230 17.455 698.395 17.835 ;
        RECT 700.870 17.455 703.035 17.835 ;
        RECT 705.510 17.455 707.675 17.835 ;
        RECT 710.150 17.455 712.315 17.835 ;
        RECT 714.790 17.455 716.955 17.835 ;
        RECT 682.335 17.175 684.450 17.455 ;
        RECT 686.975 17.175 689.090 17.455 ;
        RECT 691.615 17.175 693.730 17.455 ;
        RECT 696.255 17.175 698.370 17.455 ;
        RECT 700.895 17.175 703.010 17.455 ;
        RECT 705.535 17.175 707.650 17.455 ;
        RECT 710.175 17.175 712.290 17.455 ;
        RECT 714.815 17.175 716.930 17.455 ;
        RECT 682.310 16.795 684.475 17.175 ;
        RECT 686.950 16.795 689.115 17.175 ;
        RECT 691.590 16.795 693.755 17.175 ;
        RECT 696.230 16.795 698.395 17.175 ;
        RECT 700.870 16.795 703.035 17.175 ;
        RECT 705.510 16.795 707.675 17.175 ;
        RECT 710.150 16.795 712.315 17.175 ;
        RECT 714.790 16.795 716.955 17.175 ;
        RECT 682.335 16.515 684.450 16.795 ;
        RECT 686.975 16.515 689.090 16.795 ;
        RECT 691.615 16.515 693.730 16.795 ;
        RECT 696.255 16.515 698.370 16.795 ;
        RECT 700.895 16.515 703.010 16.795 ;
        RECT 705.535 16.515 707.650 16.795 ;
        RECT 710.175 16.515 712.290 16.795 ;
        RECT 714.815 16.515 716.930 16.795 ;
        RECT 682.310 16.135 684.475 16.515 ;
        RECT 686.950 16.135 689.115 16.515 ;
        RECT 691.590 16.135 693.755 16.515 ;
        RECT 696.230 16.135 698.395 16.515 ;
        RECT 700.870 16.135 703.035 16.515 ;
        RECT 705.510 16.135 707.675 16.515 ;
        RECT 710.150 16.135 712.315 16.515 ;
        RECT 714.790 16.135 716.955 16.515 ;
        RECT 682.335 15.855 684.450 16.135 ;
        RECT 686.975 15.855 689.090 16.135 ;
        RECT 691.615 15.855 693.730 16.135 ;
        RECT 696.255 15.855 698.370 16.135 ;
        RECT 700.895 15.855 703.010 16.135 ;
        RECT 705.535 15.855 707.650 16.135 ;
        RECT 710.175 15.855 712.290 16.135 ;
        RECT 714.815 15.855 716.930 16.135 ;
        RECT 682.310 15.475 684.475 15.855 ;
        RECT 686.950 15.475 689.115 15.855 ;
        RECT 691.590 15.475 693.755 15.855 ;
        RECT 696.230 15.475 698.395 15.855 ;
        RECT 700.870 15.475 703.035 15.855 ;
        RECT 705.510 15.475 707.675 15.855 ;
        RECT 710.150 15.475 712.315 15.855 ;
        RECT 714.790 15.475 716.955 15.855 ;
        RECT 682.335 15.195 684.450 15.475 ;
        RECT 686.975 15.195 689.090 15.475 ;
        RECT 691.615 15.195 693.730 15.475 ;
        RECT 696.255 15.195 698.370 15.475 ;
        RECT 700.895 15.195 703.010 15.475 ;
        RECT 705.535 15.195 707.650 15.475 ;
        RECT 710.175 15.195 712.290 15.475 ;
        RECT 714.815 15.195 716.930 15.475 ;
        RECT 682.310 14.815 684.475 15.195 ;
        RECT 686.950 14.815 689.115 15.195 ;
        RECT 691.590 14.815 693.755 15.195 ;
        RECT 696.230 14.815 698.395 15.195 ;
        RECT 700.870 14.815 703.035 15.195 ;
        RECT 705.510 14.815 707.675 15.195 ;
        RECT 710.150 14.815 712.315 15.195 ;
        RECT 714.790 14.815 716.955 15.195 ;
        RECT 682.335 14.535 684.450 14.815 ;
        RECT 686.975 14.535 689.090 14.815 ;
        RECT 691.615 14.535 693.730 14.815 ;
        RECT 696.255 14.535 698.370 14.815 ;
        RECT 700.895 14.535 703.010 14.815 ;
        RECT 705.535 14.535 707.650 14.815 ;
        RECT 710.175 14.535 712.290 14.815 ;
        RECT 714.815 14.535 716.930 14.815 ;
        RECT 682.310 14.155 684.475 14.535 ;
        RECT 686.950 14.155 689.115 14.535 ;
        RECT 691.590 14.155 693.755 14.535 ;
        RECT 696.230 14.155 698.395 14.535 ;
        RECT 700.870 14.155 703.035 14.535 ;
        RECT 705.510 14.155 707.675 14.535 ;
        RECT 710.150 14.155 712.315 14.535 ;
        RECT 714.790 14.155 716.955 14.535 ;
        RECT 682.335 13.875 684.450 14.155 ;
        RECT 686.975 13.875 689.090 14.155 ;
        RECT 691.615 13.875 693.730 14.155 ;
        RECT 696.255 13.875 698.370 14.155 ;
        RECT 700.895 13.875 703.010 14.155 ;
        RECT 705.535 13.875 707.650 14.155 ;
        RECT 710.175 13.875 712.290 14.155 ;
        RECT 714.815 13.875 716.930 14.155 ;
        RECT 682.310 13.495 684.475 13.875 ;
        RECT 686.950 13.495 689.115 13.875 ;
        RECT 691.590 13.495 693.755 13.875 ;
        RECT 696.230 13.495 698.395 13.875 ;
        RECT 700.870 13.495 703.035 13.875 ;
        RECT 705.510 13.495 707.675 13.875 ;
        RECT 710.150 13.495 712.315 13.875 ;
        RECT 714.790 13.495 716.955 13.875 ;
        RECT 682.335 13.215 684.450 13.495 ;
        RECT 686.975 13.215 689.090 13.495 ;
        RECT 691.615 13.215 693.730 13.495 ;
        RECT 696.255 13.215 698.370 13.495 ;
        RECT 700.895 13.215 703.010 13.495 ;
        RECT 705.535 13.215 707.650 13.495 ;
        RECT 710.175 13.215 712.290 13.495 ;
        RECT 714.815 13.215 716.930 13.495 ;
        RECT 682.310 12.835 684.475 13.215 ;
        RECT 686.950 12.835 689.115 13.215 ;
        RECT 691.590 12.835 693.755 13.215 ;
        RECT 696.230 12.835 698.395 13.215 ;
        RECT 700.870 12.835 703.035 13.215 ;
        RECT 705.510 12.835 707.675 13.215 ;
        RECT 710.150 12.835 712.315 13.215 ;
        RECT 714.790 12.835 716.955 13.215 ;
        RECT 682.335 12.555 684.450 12.835 ;
        RECT 686.975 12.555 689.090 12.835 ;
        RECT 691.615 12.555 693.730 12.835 ;
        RECT 696.255 12.555 698.370 12.835 ;
        RECT 700.895 12.555 703.010 12.835 ;
        RECT 705.535 12.555 707.650 12.835 ;
        RECT 710.175 12.555 712.290 12.835 ;
        RECT 714.815 12.555 716.930 12.835 ;
        RECT 682.310 12.175 684.475 12.555 ;
        RECT 686.950 12.175 689.115 12.555 ;
        RECT 691.590 12.175 693.755 12.555 ;
        RECT 696.230 12.175 698.395 12.555 ;
        RECT 700.870 12.175 703.035 12.555 ;
        RECT 705.510 12.175 707.675 12.555 ;
        RECT 710.150 12.175 712.315 12.555 ;
        RECT 714.790 12.175 716.955 12.555 ;
        RECT 682.335 11.895 684.450 12.175 ;
        RECT 686.975 11.895 689.090 12.175 ;
        RECT 691.615 11.895 693.730 12.175 ;
        RECT 696.255 11.895 698.370 12.175 ;
        RECT 700.895 11.895 703.010 12.175 ;
        RECT 705.535 11.895 707.650 12.175 ;
        RECT 710.175 11.895 712.290 12.175 ;
        RECT 714.815 11.895 716.930 12.175 ;
        RECT 682.310 11.515 684.475 11.895 ;
        RECT 686.950 11.515 689.115 11.895 ;
        RECT 691.590 11.515 693.755 11.895 ;
        RECT 696.230 11.515 698.395 11.895 ;
        RECT 700.870 11.515 703.035 11.895 ;
        RECT 705.510 11.515 707.675 11.895 ;
        RECT 710.150 11.515 712.315 11.895 ;
        RECT 714.790 11.515 716.955 11.895 ;
        RECT 682.335 11.235 684.450 11.515 ;
        RECT 686.975 11.235 689.090 11.515 ;
        RECT 691.615 11.235 693.730 11.515 ;
        RECT 696.255 11.235 698.370 11.515 ;
        RECT 700.895 11.235 703.010 11.515 ;
        RECT 705.535 11.235 707.650 11.515 ;
        RECT 710.175 11.235 712.290 11.515 ;
        RECT 714.815 11.235 716.930 11.515 ;
        RECT 682.310 10.855 684.475 11.235 ;
        RECT 686.950 10.855 689.115 11.235 ;
        RECT 691.590 10.855 693.755 11.235 ;
        RECT 696.230 10.855 698.395 11.235 ;
        RECT 700.870 10.855 703.035 11.235 ;
        RECT 705.510 10.855 707.675 11.235 ;
        RECT 710.150 10.855 712.315 11.235 ;
        RECT 714.790 10.855 716.955 11.235 ;
        RECT 682.335 10.575 684.450 10.855 ;
        RECT 686.975 10.575 689.090 10.855 ;
        RECT 691.615 10.575 693.730 10.855 ;
        RECT 696.255 10.575 698.370 10.855 ;
        RECT 700.895 10.575 703.010 10.855 ;
        RECT 705.535 10.575 707.650 10.855 ;
        RECT 710.175 10.575 712.290 10.855 ;
        RECT 714.815 10.575 716.930 10.855 ;
        RECT 682.310 10.195 684.475 10.575 ;
        RECT 686.950 10.195 689.115 10.575 ;
        RECT 691.590 10.195 693.755 10.575 ;
        RECT 696.230 10.195 698.395 10.575 ;
        RECT 700.870 10.195 703.035 10.575 ;
        RECT 705.510 10.195 707.675 10.575 ;
        RECT 710.150 10.195 712.315 10.575 ;
        RECT 714.790 10.195 716.955 10.575 ;
        RECT 682.335 9.915 684.450 10.195 ;
        RECT 686.975 9.915 689.090 10.195 ;
        RECT 691.615 9.915 693.730 10.195 ;
        RECT 696.255 9.915 698.370 10.195 ;
        RECT 700.895 9.915 703.010 10.195 ;
        RECT 705.535 9.915 707.650 10.195 ;
        RECT 710.175 9.915 712.290 10.195 ;
        RECT 714.815 9.915 716.930 10.195 ;
        RECT 682.310 9.535 684.475 9.915 ;
        RECT 686.950 9.535 689.115 9.915 ;
        RECT 691.590 9.535 693.755 9.915 ;
        RECT 696.230 9.535 698.395 9.915 ;
        RECT 700.870 9.535 703.035 9.915 ;
        RECT 705.510 9.535 707.675 9.915 ;
        RECT 710.150 9.535 712.315 9.915 ;
        RECT 714.790 9.535 716.955 9.915 ;
        RECT 682.335 9.255 684.450 9.535 ;
        RECT 686.975 9.255 689.090 9.535 ;
        RECT 691.615 9.255 693.730 9.535 ;
        RECT 696.255 9.255 698.370 9.535 ;
        RECT 700.895 9.255 703.010 9.535 ;
        RECT 705.535 9.255 707.650 9.535 ;
        RECT 710.175 9.255 712.290 9.535 ;
        RECT 714.815 9.255 716.930 9.535 ;
        RECT 682.310 8.875 684.475 9.255 ;
        RECT 686.950 8.875 689.115 9.255 ;
        RECT 691.590 8.875 693.755 9.255 ;
        RECT 696.230 8.875 698.395 9.255 ;
        RECT 700.870 8.875 703.035 9.255 ;
        RECT 705.510 8.875 707.675 9.255 ;
        RECT 710.150 8.875 712.315 9.255 ;
        RECT 714.790 8.875 716.955 9.255 ;
        RECT 682.335 2.500 684.450 8.875 ;
        RECT 686.975 2.500 689.090 8.875 ;
        RECT 691.615 2.500 693.730 8.875 ;
        RECT 696.255 2.500 698.370 8.875 ;
        RECT 700.895 2.500 703.010 8.875 ;
        RECT 705.535 2.500 707.650 8.875 ;
        RECT 710.175 2.500 712.290 8.875 ;
        RECT 714.815 2.500 716.930 8.875 ;
        RECT 0.000 0.000 717.540 2.500 ;
    END
  END VDD
  OBS
      LAYER Metal1 ;
              RECT 3.905 11.185 8.285 17.775 ;
        RECT 14.281 11.185 18.661 17.775 ;
        RECT 24.657 11.185 29.037 17.775 ;
        RECT 35.033 11.185 39.413 17.775 ;
        RECT 46.409 11.185 50.789 17.775 ;
        RECT 56.785 11.185 61.165 17.775 ;
        RECT 67.161 11.185 71.541 17.775 ;
        RECT 77.537 11.185 81.917 17.775 ;
        RECT 88.913 11.185 93.293 17.775 ;
        RECT 99.289 11.185 103.669 17.775 ;
        RECT 109.665 11.185 114.045 17.775 ;
        RECT 120.041 11.185 124.421 17.775 ;
        RECT 131.417 11.185 135.797 17.775 ;
        RECT 141.793 11.185 146.173 17.775 ;
        RECT 152.169 11.185 156.549 17.775 ;
        RECT 162.545 11.185 166.925 17.775 ;
        RECT 173.921 11.185 178.301 17.775 ;
        RECT 184.297 11.185 188.677 17.775 ;
        RECT 194.673 11.185 199.053 17.775 ;
        RECT 205.049 11.185 209.429 17.775 ;
        RECT 216.425 11.185 220.805 17.775 ;
        RECT 226.801 11.185 231.181 17.775 ;
        RECT 237.177 11.185 241.557 17.775 ;
        RECT 247.553 11.185 251.933 17.775 ;
        RECT 258.929 11.185 263.309 17.775 ;
        RECT 269.305 11.185 273.685 17.775 ;
        RECT 279.681 11.185 284.061 17.775 ;
        RECT 290.057 11.185 294.437 17.775 ;
        RECT 301.433 11.185 305.813 17.775 ;
        RECT 311.809 11.185 316.189 17.775 ;
        RECT 322.185 11.185 326.565 17.775 ;
        RECT 332.561 11.185 336.941 17.775 ;
        RECT 343.937 11.185 348.317 17.775 ;
        RECT 354.313 11.185 358.693 17.775 ;
        RECT 364.689 11.185 369.069 17.775 ;
        RECT 375.065 11.185 379.445 17.775 ;
        RECT 386.441 11.185 390.821 17.775 ;
        RECT 396.817 11.185 401.197 17.775 ;
        RECT 407.193 11.185 411.573 17.775 ;
        RECT 417.569 11.185 421.949 17.775 ;
        RECT 428.945 11.185 433.325 17.775 ;
        RECT 439.321 11.185 443.701 17.775 ;
        RECT 449.697 11.185 454.077 17.775 ;
        RECT 460.073 11.185 464.453 17.775 ;
        RECT 471.449 11.185 475.829 17.775 ;
        RECT 481.825 11.185 486.205 17.775 ;
        RECT 492.201 11.185 496.581 17.775 ;
        RECT 502.577 11.185 506.957 17.775 ;
        RECT 513.953 11.185 518.333 17.775 ;
        RECT 524.329 11.185 528.709 17.775 ;
        RECT 534.705 11.185 539.085 17.775 ;
        RECT 545.081 11.185 549.461 17.775 ;
        RECT 556.457 11.185 560.837 17.775 ;
        RECT 566.833 11.185 571.213 17.775 ;
        RECT 577.209 11.185 581.589 17.775 ;
        RECT 587.585 11.185 591.965 17.775 ;
        RECT 598.961 11.185 603.341 17.775 ;
        RECT 609.337 11.185 613.717 17.775 ;
        RECT 619.713 11.185 624.093 17.775 ;
        RECT 630.089 11.185 634.469 17.775 ;
        RECT 641.465 11.185 645.845 17.775 ;
        RECT 651.841 11.185 656.221 17.775 ;
        RECT 662.217 11.185 666.597 17.775 ;
        RECT 672.593 11.185 676.973 17.775 ;
        RECT 3.915 49.781 8.295 56.371 ;
        RECT 14.291 49.781 18.671 56.371 ;
        RECT 24.667 49.781 29.047 56.371 ;
        RECT 35.043 49.781 39.423 56.371 ;
        RECT 46.419 49.781 50.799 56.371 ;
        RECT 56.795 49.781 61.175 56.371 ;
        RECT 67.171 49.781 71.551 56.371 ;
        RECT 77.547 49.781 81.927 56.371 ;
        RECT 88.923 49.781 93.303 56.371 ;
        RECT 99.299 49.781 103.679 56.371 ;
        RECT 109.675 49.781 114.055 56.371 ;
        RECT 120.051 49.781 124.431 56.371 ;
        RECT 131.427 49.781 135.807 56.371 ;
        RECT 141.803 49.781 146.183 56.371 ;
        RECT 152.179 49.781 156.559 56.371 ;
        RECT 162.555 49.781 166.935 56.371 ;
        RECT 173.931 49.781 178.311 56.371 ;
        RECT 184.307 49.781 188.687 56.371 ;
        RECT 194.683 49.781 199.063 56.371 ;
        RECT 205.059 49.781 209.439 56.371 ;
        RECT 216.435 49.781 220.815 56.371 ;
        RECT 226.811 49.781 231.191 56.371 ;
        RECT 237.187 49.781 241.567 56.371 ;
        RECT 247.563 49.781 251.943 56.371 ;
        RECT 258.939 49.781 263.319 56.371 ;
        RECT 269.315 49.781 273.695 56.371 ;
        RECT 279.691 49.781 284.071 56.371 ;
        RECT 290.067 49.781 294.447 56.371 ;
        RECT 301.443 49.781 305.823 56.371 ;
        RECT 311.819 49.781 316.199 56.371 ;
        RECT 322.195 49.781 326.575 56.371 ;
        RECT 332.571 49.781 336.951 56.371 ;
        RECT 343.947 49.781 348.327 56.371 ;
        RECT 354.323 49.781 358.703 56.371 ;
        RECT 364.699 49.781 369.079 56.371 ;
        RECT 375.075 49.781 379.455 56.371 ;
        RECT 386.451 49.781 390.831 56.371 ;
        RECT 396.827 49.781 401.207 56.371 ;
        RECT 407.203 49.781 411.583 56.371 ;
        RECT 417.579 49.781 421.959 56.371 ;
        RECT 428.955 49.781 433.335 56.371 ;
        RECT 439.331 49.781 443.711 56.371 ;
        RECT 449.707 49.781 454.087 56.371 ;
        RECT 460.083 49.781 464.463 56.371 ;
        RECT 471.459 49.781 475.839 56.371 ;
        RECT 481.835 49.781 486.215 56.371 ;
        RECT 492.211 49.781 496.591 56.371 ;
        RECT 502.587 49.781 506.967 56.371 ;
        RECT 513.963 49.781 518.343 56.371 ;
        RECT 524.339 49.781 528.719 56.371 ;
        RECT 534.715 49.781 539.095 56.371 ;
        RECT 545.091 49.781 549.471 56.371 ;
        RECT 556.467 49.781 560.847 56.371 ;
        RECT 566.843 49.781 571.223 56.371 ;
        RECT 577.219 49.781 581.599 56.371 ;
        RECT 587.595 49.781 591.975 56.371 ;
        RECT 598.971 49.781 603.351 56.371 ;
        RECT 609.347 49.781 613.727 56.371 ;
        RECT 619.723 49.781 624.103 56.371 ;
        RECT 630.099 49.781 634.479 56.371 ;
        RECT 641.475 49.781 645.855 56.371 ;
        RECT 651.851 49.781 656.231 56.371 ;
        RECT 662.227 49.781 666.607 56.371 ;
        RECT 672.603 49.781 676.983 56.371 ;

        RECT 1.975 59.605 2.675 60.305 ;
        RECT 0.735 9.370 1.905 59.380 ;
        RECT 1.525 9.360 1.905 9.370 ;
        RECT 2.755 56.865 6.970 59.380 ;
        RECT 2.755 9.360 3.125 56.865 ;
        RECT 5.220 54.845 6.970 56.865 ;
        RECT 5.690 49.385 6.500 53.395 ;
        RECT 5.250 46.485 6.950 49.385 ;
        RECT 5.250 19.685 6.950 22.585 ;
        RECT 5.700 15.660 6.510 19.685 ;
        RECT 5.230 12.190 6.980 14.210 ;
        RECT 9.075 12.190 9.445 59.695 ;
        RECT 5.230 9.675 9.445 12.190 ;
        RECT 10.295 59.685 10.675 59.695 ;
        RECT 11.815 59.685 12.195 59.695 ;
        RECT 10.295 9.675 12.195 59.685 ;
        RECT 13.045 12.190 13.415 59.695 ;
        RECT 19.810 59.605 20.510 60.305 ;
        RECT 22.550 59.605 23.250 60.305 ;
        RECT 15.515 56.865 19.730 59.380 ;
        RECT 15.515 54.845 17.265 56.865 ;
        RECT 15.985 49.385 16.795 53.395 ;
        RECT 15.550 43.785 17.250 49.385 ;
        RECT 15.550 19.685 17.250 25.285 ;
        RECT 15.980 15.660 16.790 19.685 ;
        RECT 15.510 12.190 17.260 14.210 ;
        RECT 13.045 9.675 17.260 12.190 ;
        RECT 9.525 8.750 10.225 9.450 ;
        RECT 12.265 8.750 12.965 9.450 ;
        RECT 19.360 9.360 19.730 56.865 ;
        RECT 20.580 9.370 22.480 59.380 ;
        RECT 20.580 9.360 20.960 9.370 ;
        RECT 22.100 9.360 22.480 9.370 ;
        RECT 23.330 56.865 27.545 59.380 ;
        RECT 23.330 9.360 23.700 56.865 ;
        RECT 25.795 54.845 27.545 56.865 ;
        RECT 26.265 49.385 27.075 53.395 ;
        RECT 25.825 41.085 27.525 49.385 ;
        RECT 25.825 19.685 27.525 27.985 ;
        RECT 26.275 15.660 27.085 19.685 ;
        RECT 25.805 12.190 27.555 14.210 ;
        RECT 29.650 12.190 30.020 59.695 ;
        RECT 25.805 9.675 30.020 12.190 ;
        RECT 30.870 59.685 31.250 59.695 ;
        RECT 32.390 59.685 32.770 59.695 ;
        RECT 30.870 9.675 32.770 59.685 ;
        RECT 33.620 12.190 33.990 59.695 ;
        RECT 40.385 59.605 41.085 60.305 ;
        RECT 44.545 59.605 45.245 60.305 ;
        RECT 36.090 56.865 40.305 59.380 ;
        RECT 36.090 54.845 37.840 56.865 ;
        RECT 36.560 49.385 37.370 53.395 ;
        RECT 36.125 38.385 37.825 49.385 ;
        RECT 36.125 19.685 37.825 30.685 ;
        RECT 36.555 15.660 37.365 19.685 ;
        RECT 36.085 12.190 37.835 14.210 ;
        RECT 33.620 9.675 37.835 12.190 ;
        RECT 30.100 8.750 30.800 9.450 ;
        RECT 32.840 8.750 33.540 9.450 ;
        RECT 39.935 9.360 40.305 56.865 ;
        RECT 41.155 9.370 42.325 59.380 ;
        RECT 43.305 9.370 44.475 59.380 ;
        RECT 41.155 9.360 41.535 9.370 ;
        RECT 44.095 9.360 44.475 9.370 ;
        RECT 45.325 56.865 49.540 59.380 ;
        RECT 45.325 9.360 45.695 56.865 ;
        RECT 47.790 54.845 49.540 56.865 ;
        RECT 48.260 49.385 49.070 53.395 ;
        RECT 47.820 46.485 49.520 49.385 ;
        RECT 47.820 19.685 49.520 22.585 ;
        RECT 48.270 15.660 49.080 19.685 ;
        RECT 47.800 12.190 49.550 14.210 ;
        RECT 51.645 12.190 52.015 59.695 ;
        RECT 47.800 9.675 52.015 12.190 ;
        RECT 52.865 59.685 53.245 59.695 ;
        RECT 54.385 59.685 54.765 59.695 ;
        RECT 52.865 9.675 54.765 59.685 ;
        RECT 55.615 12.190 55.985 59.695 ;
        RECT 62.380 59.605 63.080 60.305 ;
        RECT 65.120 59.605 65.820 60.305 ;
        RECT 58.085 56.865 62.300 59.380 ;
        RECT 58.085 54.845 59.835 56.865 ;
        RECT 58.555 49.385 59.365 53.395 ;
        RECT 58.120 43.785 59.820 49.385 ;
        RECT 58.120 19.685 59.820 25.285 ;
        RECT 58.550 15.660 59.360 19.685 ;
        RECT 58.080 12.190 59.830 14.210 ;
        RECT 55.615 9.675 59.830 12.190 ;
        RECT 52.095 8.750 52.795 9.450 ;
        RECT 54.835 8.750 55.535 9.450 ;
        RECT 61.930 9.360 62.300 56.865 ;
        RECT 63.150 9.370 65.050 59.380 ;
        RECT 63.150 9.360 63.530 9.370 ;
        RECT 64.670 9.360 65.050 9.370 ;
        RECT 65.900 56.865 70.115 59.380 ;
        RECT 65.900 9.360 66.270 56.865 ;
        RECT 68.365 54.845 70.115 56.865 ;
        RECT 68.835 49.385 69.645 53.395 ;
        RECT 68.395 41.085 70.095 49.385 ;
        RECT 68.395 19.685 70.095 27.985 ;
        RECT 68.845 15.660 69.655 19.685 ;
        RECT 68.375 12.190 70.125 14.210 ;
        RECT 72.220 12.190 72.590 59.695 ;
        RECT 68.375 9.675 72.590 12.190 ;
        RECT 73.440 59.685 73.820 59.695 ;
        RECT 74.960 59.685 75.340 59.695 ;
        RECT 73.440 9.675 75.340 59.685 ;
        RECT 76.190 12.190 76.560 59.695 ;
        RECT 82.955 59.605 83.655 60.305 ;
        RECT 87.115 59.605 87.815 60.305 ;
        RECT 78.660 56.865 82.875 59.380 ;
        RECT 78.660 54.845 80.410 56.865 ;
        RECT 79.130 49.385 79.940 53.395 ;
        RECT 78.695 38.385 80.395 49.385 ;
        RECT 78.695 19.685 80.395 30.685 ;
        RECT 79.125 15.660 79.935 19.685 ;
        RECT 78.655 12.190 80.405 14.210 ;
        RECT 76.190 9.675 80.405 12.190 ;
        RECT 72.670 8.750 73.370 9.450 ;
        RECT 75.410 8.750 76.110 9.450 ;
        RECT 82.505 9.360 82.875 56.865 ;
        RECT 83.725 9.370 84.895 59.380 ;
        RECT 85.875 9.370 87.045 59.380 ;
        RECT 83.725 9.360 84.105 9.370 ;
        RECT 86.665 9.360 87.045 9.370 ;
        RECT 87.895 56.865 92.110 59.380 ;
        RECT 87.895 9.360 88.265 56.865 ;
        RECT 90.360 54.845 92.110 56.865 ;
        RECT 90.830 49.385 91.640 53.395 ;
        RECT 90.390 46.485 92.090 49.385 ;
        RECT 90.390 19.685 92.090 22.585 ;
        RECT 90.840 15.660 91.650 19.685 ;
        RECT 90.370 12.190 92.120 14.210 ;
        RECT 94.215 12.190 94.585 59.695 ;
        RECT 90.370 9.675 94.585 12.190 ;
        RECT 95.435 59.685 95.815 59.695 ;
        RECT 96.955 59.685 97.335 59.695 ;
        RECT 95.435 9.675 97.335 59.685 ;
        RECT 98.185 12.190 98.555 59.695 ;
        RECT 104.950 59.605 105.650 60.305 ;
        RECT 107.690 59.605 108.390 60.305 ;
        RECT 100.655 56.865 104.870 59.380 ;
        RECT 100.655 54.845 102.405 56.865 ;
        RECT 101.125 49.385 101.935 53.395 ;
        RECT 100.690 43.785 102.390 49.385 ;
        RECT 100.690 19.685 102.390 25.285 ;
        RECT 101.120 15.660 101.930 19.685 ;
        RECT 100.650 12.190 102.400 14.210 ;
        RECT 98.185 9.675 102.400 12.190 ;
        RECT 94.665 8.750 95.365 9.450 ;
        RECT 97.405 8.750 98.105 9.450 ;
        RECT 104.500 9.360 104.870 56.865 ;
        RECT 105.720 9.370 107.620 59.380 ;
        RECT 105.720 9.360 106.100 9.370 ;
        RECT 107.240 9.360 107.620 9.370 ;
        RECT 108.470 56.865 112.685 59.380 ;
        RECT 108.470 9.360 108.840 56.865 ;
        RECT 110.935 54.845 112.685 56.865 ;
        RECT 111.405 49.385 112.215 53.395 ;
        RECT 110.965 41.085 112.665 49.385 ;
        RECT 110.965 19.685 112.665 27.985 ;
        RECT 111.415 15.660 112.225 19.685 ;
        RECT 110.945 12.190 112.695 14.210 ;
        RECT 114.790 12.190 115.160 59.695 ;
        RECT 110.945 9.675 115.160 12.190 ;
        RECT 116.010 59.685 116.390 59.695 ;
        RECT 117.530 59.685 117.910 59.695 ;
        RECT 116.010 9.675 117.910 59.685 ;
        RECT 118.760 12.190 119.130 59.695 ;
        RECT 125.525 59.605 126.225 60.305 ;
        RECT 129.685 59.605 130.385 60.305 ;
        RECT 121.230 56.865 125.445 59.380 ;
        RECT 121.230 54.845 122.980 56.865 ;
        RECT 121.700 49.385 122.510 53.395 ;
        RECT 121.265 38.385 122.965 49.385 ;
        RECT 121.265 19.685 122.965 30.685 ;
        RECT 121.695 15.660 122.505 19.685 ;
        RECT 121.225 12.190 122.975 14.210 ;
        RECT 118.760 9.675 122.975 12.190 ;
        RECT 115.240 8.750 115.940 9.450 ;
        RECT 117.980 8.750 118.680 9.450 ;
        RECT 125.075 9.360 125.445 56.865 ;
        RECT 126.295 9.370 127.465 59.380 ;
        RECT 128.445 9.370 129.615 59.380 ;
        RECT 126.295 9.360 126.675 9.370 ;
        RECT 129.235 9.360 129.615 9.370 ;
        RECT 130.465 56.865 134.680 59.380 ;
        RECT 130.465 9.360 130.835 56.865 ;
        RECT 132.930 54.845 134.680 56.865 ;
        RECT 133.400 49.385 134.210 53.395 ;
        RECT 132.960 46.485 134.660 49.385 ;
        RECT 132.960 19.685 134.660 22.585 ;
        RECT 133.410 15.660 134.220 19.685 ;
        RECT 132.940 12.190 134.690 14.210 ;
        RECT 136.785 12.190 137.155 59.695 ;
        RECT 132.940 9.675 137.155 12.190 ;
        RECT 138.005 59.685 138.385 59.695 ;
        RECT 139.525 59.685 139.905 59.695 ;
        RECT 138.005 9.675 139.905 59.685 ;
        RECT 140.755 12.190 141.125 59.695 ;
        RECT 147.520 59.605 148.220 60.305 ;
        RECT 150.260 59.605 150.960 60.305 ;
        RECT 143.225 56.865 147.440 59.380 ;
        RECT 143.225 54.845 144.975 56.865 ;
        RECT 143.695 49.385 144.505 53.395 ;
        RECT 143.260 43.785 144.960 49.385 ;
        RECT 143.260 19.685 144.960 25.285 ;
        RECT 143.690 15.660 144.500 19.685 ;
        RECT 143.220 12.190 144.970 14.210 ;
        RECT 140.755 9.675 144.970 12.190 ;
        RECT 137.235 8.750 137.935 9.450 ;
        RECT 139.975 8.750 140.675 9.450 ;
        RECT 147.070 9.360 147.440 56.865 ;
        RECT 148.290 9.370 150.190 59.380 ;
        RECT 148.290 9.360 148.670 9.370 ;
        RECT 149.810 9.360 150.190 9.370 ;
        RECT 151.040 56.865 155.255 59.380 ;
        RECT 151.040 9.360 151.410 56.865 ;
        RECT 153.505 54.845 155.255 56.865 ;
        RECT 153.975 49.385 154.785 53.395 ;
        RECT 153.535 41.085 155.235 49.385 ;
        RECT 153.535 19.685 155.235 27.985 ;
        RECT 153.985 15.660 154.795 19.685 ;
        RECT 153.515 12.190 155.265 14.210 ;
        RECT 157.360 12.190 157.730 59.695 ;
        RECT 153.515 9.675 157.730 12.190 ;
        RECT 158.580 59.685 158.960 59.695 ;
        RECT 160.100 59.685 160.480 59.695 ;
        RECT 158.580 9.675 160.480 59.685 ;
        RECT 161.330 12.190 161.700 59.695 ;
        RECT 168.095 59.605 168.795 60.305 ;
        RECT 172.255 59.605 172.955 60.305 ;
        RECT 163.800 56.865 168.015 59.380 ;
        RECT 163.800 54.845 165.550 56.865 ;
        RECT 164.270 49.385 165.080 53.395 ;
        RECT 163.835 38.385 165.535 49.385 ;
        RECT 163.835 19.685 165.535 30.685 ;
        RECT 164.265 15.660 165.075 19.685 ;
        RECT 163.795 12.190 165.545 14.210 ;
        RECT 161.330 9.675 165.545 12.190 ;
        RECT 157.810 8.750 158.510 9.450 ;
        RECT 160.550 8.750 161.250 9.450 ;
        RECT 167.645 9.360 168.015 56.865 ;
        RECT 168.865 9.370 170.035 59.380 ;
        RECT 171.015 9.370 172.185 59.380 ;
        RECT 168.865 9.360 169.245 9.370 ;
        RECT 171.805 9.360 172.185 9.370 ;
        RECT 173.035 56.865 177.250 59.380 ;
        RECT 173.035 9.360 173.405 56.865 ;
        RECT 175.500 54.845 177.250 56.865 ;
        RECT 175.970 49.385 176.780 53.395 ;
        RECT 175.530 46.485 177.230 49.385 ;
        RECT 175.530 19.685 177.230 22.585 ;
        RECT 175.980 15.660 176.790 19.685 ;
        RECT 175.510 12.190 177.260 14.210 ;
        RECT 179.355 12.190 179.725 59.695 ;
        RECT 175.510 9.675 179.725 12.190 ;
        RECT 180.575 59.685 180.955 59.695 ;
        RECT 182.095 59.685 182.475 59.695 ;
        RECT 180.575 9.675 182.475 59.685 ;
        RECT 183.325 12.190 183.695 59.695 ;
        RECT 190.090 59.605 190.790 60.305 ;
        RECT 192.830 59.605 193.530 60.305 ;
        RECT 185.795 56.865 190.010 59.380 ;
        RECT 185.795 54.845 187.545 56.865 ;
        RECT 186.265 49.385 187.075 53.395 ;
        RECT 185.830 43.785 187.530 49.385 ;
        RECT 185.830 19.685 187.530 25.285 ;
        RECT 186.260 15.660 187.070 19.685 ;
        RECT 185.790 12.190 187.540 14.210 ;
        RECT 183.325 9.675 187.540 12.190 ;
        RECT 179.805 8.750 180.505 9.450 ;
        RECT 182.545 8.750 183.245 9.450 ;
        RECT 189.640 9.360 190.010 56.865 ;
        RECT 190.860 9.370 192.760 59.380 ;
        RECT 190.860 9.360 191.240 9.370 ;
        RECT 192.380 9.360 192.760 9.370 ;
        RECT 193.610 56.865 197.825 59.380 ;
        RECT 193.610 9.360 193.980 56.865 ;
        RECT 196.075 54.845 197.825 56.865 ;
        RECT 196.545 49.385 197.355 53.395 ;
        RECT 196.105 41.085 197.805 49.385 ;
        RECT 196.105 19.685 197.805 27.985 ;
        RECT 196.555 15.660 197.365 19.685 ;
        RECT 196.085 12.190 197.835 14.210 ;
        RECT 199.930 12.190 200.300 59.695 ;
        RECT 196.085 9.675 200.300 12.190 ;
        RECT 201.150 59.685 201.530 59.695 ;
        RECT 202.670 59.685 203.050 59.695 ;
        RECT 201.150 9.675 203.050 59.685 ;
        RECT 203.900 12.190 204.270 59.695 ;
        RECT 210.665 59.605 211.365 60.305 ;
        RECT 214.825 59.605 215.525 60.305 ;
        RECT 206.370 56.865 210.585 59.380 ;
        RECT 206.370 54.845 208.120 56.865 ;
        RECT 206.840 49.385 207.650 53.395 ;
        RECT 206.405 38.385 208.105 49.385 ;
        RECT 206.405 19.685 208.105 30.685 ;
        RECT 206.835 15.660 207.645 19.685 ;
        RECT 206.365 12.190 208.115 14.210 ;
        RECT 203.900 9.675 208.115 12.190 ;
        RECT 200.380 8.750 201.080 9.450 ;
        RECT 203.120 8.750 203.820 9.450 ;
        RECT 210.215 9.360 210.585 56.865 ;
        RECT 211.435 9.370 212.605 59.380 ;
        RECT 213.585 9.370 214.755 59.380 ;
        RECT 211.435 9.360 211.815 9.370 ;
        RECT 214.375 9.360 214.755 9.370 ;
        RECT 215.605 56.865 219.820 59.380 ;
        RECT 215.605 9.360 215.975 56.865 ;
        RECT 218.070 54.845 219.820 56.865 ;
        RECT 218.540 49.385 219.350 53.395 ;
        RECT 218.100 46.485 219.800 49.385 ;
        RECT 218.100 19.685 219.800 22.585 ;
        RECT 218.550 15.660 219.360 19.685 ;
        RECT 218.080 12.190 219.830 14.210 ;
        RECT 221.925 12.190 222.295 59.695 ;
        RECT 218.080 9.675 222.295 12.190 ;
        RECT 223.145 59.685 223.525 59.695 ;
        RECT 224.665 59.685 225.045 59.695 ;
        RECT 223.145 9.675 225.045 59.685 ;
        RECT 225.895 12.190 226.265 59.695 ;
        RECT 232.660 59.605 233.360 60.305 ;
        RECT 235.400 59.605 236.100 60.305 ;
        RECT 228.365 56.865 232.580 59.380 ;
        RECT 228.365 54.845 230.115 56.865 ;
        RECT 228.835 49.385 229.645 53.395 ;
        RECT 228.400 43.785 230.100 49.385 ;
        RECT 228.400 19.685 230.100 25.285 ;
        RECT 228.830 15.660 229.640 19.685 ;
        RECT 228.360 12.190 230.110 14.210 ;
        RECT 225.895 9.675 230.110 12.190 ;
        RECT 222.375 8.750 223.075 9.450 ;
        RECT 225.115 8.750 225.815 9.450 ;
        RECT 232.210 9.360 232.580 56.865 ;
        RECT 233.430 9.370 235.330 59.380 ;
        RECT 233.430 9.360 233.810 9.370 ;
        RECT 234.950 9.360 235.330 9.370 ;
        RECT 236.180 56.865 240.395 59.380 ;
        RECT 236.180 9.360 236.550 56.865 ;
        RECT 238.645 54.845 240.395 56.865 ;
        RECT 239.115 49.385 239.925 53.395 ;
        RECT 238.675 41.085 240.375 49.385 ;
        RECT 238.675 19.685 240.375 27.985 ;
        RECT 239.125 15.660 239.935 19.685 ;
        RECT 238.655 12.190 240.405 14.210 ;
        RECT 242.500 12.190 242.870 59.695 ;
        RECT 238.655 9.675 242.870 12.190 ;
        RECT 243.720 59.685 244.100 59.695 ;
        RECT 245.240 59.685 245.620 59.695 ;
        RECT 243.720 9.675 245.620 59.685 ;
        RECT 246.470 12.190 246.840 59.695 ;
        RECT 253.235 59.605 253.935 60.305 ;
        RECT 257.395 59.605 258.095 60.305 ;
        RECT 248.940 56.865 253.155 59.380 ;
        RECT 248.940 54.845 250.690 56.865 ;
        RECT 249.410 49.385 250.220 53.395 ;
        RECT 248.975 38.385 250.675 49.385 ;
        RECT 248.975 19.685 250.675 30.685 ;
        RECT 249.405 15.660 250.215 19.685 ;
        RECT 248.935 12.190 250.685 14.210 ;
        RECT 246.470 9.675 250.685 12.190 ;
        RECT 242.950 8.750 243.650 9.450 ;
        RECT 245.690 8.750 246.390 9.450 ;
        RECT 252.785 9.360 253.155 56.865 ;
        RECT 254.005 9.370 255.175 59.380 ;
        RECT 256.155 9.370 257.325 59.380 ;
        RECT 254.005 9.360 254.385 9.370 ;
        RECT 256.945 9.360 257.325 9.370 ;
        RECT 258.175 56.865 262.390 59.380 ;
        RECT 258.175 9.360 258.545 56.865 ;
        RECT 260.640 54.845 262.390 56.865 ;
        RECT 261.110 49.385 261.920 53.395 ;
        RECT 260.670 46.485 262.370 49.385 ;
        RECT 260.670 19.685 262.370 22.585 ;
        RECT 261.120 15.660 261.930 19.685 ;
        RECT 260.650 12.190 262.400 14.210 ;
        RECT 264.495 12.190 264.865 59.695 ;
        RECT 260.650 9.675 264.865 12.190 ;
        RECT 265.715 59.685 266.095 59.695 ;
        RECT 267.235 59.685 267.615 59.695 ;
        RECT 265.715 9.675 267.615 59.685 ;
        RECT 268.465 12.190 268.835 59.695 ;
        RECT 275.230 59.605 275.930 60.305 ;
        RECT 277.970 59.605 278.670 60.305 ;
        RECT 270.935 56.865 275.150 59.380 ;
        RECT 270.935 54.845 272.685 56.865 ;
        RECT 271.405 49.385 272.215 53.395 ;
        RECT 270.970 43.785 272.670 49.385 ;
        RECT 270.970 19.685 272.670 25.285 ;
        RECT 271.400 15.660 272.210 19.685 ;
        RECT 270.930 12.190 272.680 14.210 ;
        RECT 268.465 9.675 272.680 12.190 ;
        RECT 264.945 8.750 265.645 9.450 ;
        RECT 267.685 8.750 268.385 9.450 ;
        RECT 274.780 9.360 275.150 56.865 ;
        RECT 276.000 9.370 277.900 59.380 ;
        RECT 276.000 9.360 276.380 9.370 ;
        RECT 277.520 9.360 277.900 9.370 ;
        RECT 278.750 56.865 282.965 59.380 ;
        RECT 278.750 9.360 279.120 56.865 ;
        RECT 281.215 54.845 282.965 56.865 ;
        RECT 281.685 49.385 282.495 53.395 ;
        RECT 281.245 41.085 282.945 49.385 ;
        RECT 281.245 19.685 282.945 27.985 ;
        RECT 281.695 15.660 282.505 19.685 ;
        RECT 281.225 12.190 282.975 14.210 ;
        RECT 285.070 12.190 285.440 59.695 ;
        RECT 281.225 9.675 285.440 12.190 ;
        RECT 286.290 59.685 286.670 59.695 ;
        RECT 287.810 59.685 288.190 59.695 ;
        RECT 286.290 9.675 288.190 59.685 ;
        RECT 289.040 12.190 289.410 59.695 ;
        RECT 295.805 59.605 296.505 60.305 ;
        RECT 299.965 59.605 300.665 60.305 ;
        RECT 291.510 56.865 295.725 59.380 ;
        RECT 291.510 54.845 293.260 56.865 ;
        RECT 291.980 49.385 292.790 53.395 ;
        RECT 291.545 38.385 293.245 49.385 ;
        RECT 291.545 19.685 293.245 30.685 ;
        RECT 291.975 15.660 292.785 19.685 ;
        RECT 291.505 12.190 293.255 14.210 ;
        RECT 289.040 9.675 293.255 12.190 ;
        RECT 285.520 8.750 286.220 9.450 ;
        RECT 288.260 8.750 288.960 9.450 ;
        RECT 295.355 9.360 295.725 56.865 ;
        RECT 296.575 9.370 297.745 59.380 ;
        RECT 298.725 9.370 299.895 59.380 ;
        RECT 296.575 9.360 296.955 9.370 ;
        RECT 299.515 9.360 299.895 9.370 ;
        RECT 300.745 56.865 304.960 59.380 ;
        RECT 300.745 9.360 301.115 56.865 ;
        RECT 303.210 54.845 304.960 56.865 ;
        RECT 303.680 49.385 304.490 53.395 ;
        RECT 303.240 46.485 304.940 49.385 ;
        RECT 303.240 19.685 304.940 22.585 ;
        RECT 303.690 15.660 304.500 19.685 ;
        RECT 303.220 12.190 304.970 14.210 ;
        RECT 307.065 12.190 307.435 59.695 ;
        RECT 303.220 9.675 307.435 12.190 ;
        RECT 308.285 59.685 308.665 59.695 ;
        RECT 309.805 59.685 310.185 59.695 ;
        RECT 308.285 9.675 310.185 59.685 ;
        RECT 311.035 12.190 311.405 59.695 ;
        RECT 317.800 59.605 318.500 60.305 ;
        RECT 320.540 59.605 321.240 60.305 ;
        RECT 313.505 56.865 317.720 59.380 ;
        RECT 313.505 54.845 315.255 56.865 ;
        RECT 313.975 49.385 314.785 53.395 ;
        RECT 313.540 43.785 315.240 49.385 ;
        RECT 313.540 19.685 315.240 25.285 ;
        RECT 313.970 15.660 314.780 19.685 ;
        RECT 313.500 12.190 315.250 14.210 ;
        RECT 311.035 9.675 315.250 12.190 ;
        RECT 307.515 8.750 308.215 9.450 ;
        RECT 310.255 8.750 310.955 9.450 ;
        RECT 317.350 9.360 317.720 56.865 ;
        RECT 318.570 9.370 320.470 59.380 ;
        RECT 318.570 9.360 318.950 9.370 ;
        RECT 320.090 9.360 320.470 9.370 ;
        RECT 321.320 56.865 325.535 59.380 ;
        RECT 321.320 9.360 321.690 56.865 ;
        RECT 323.785 54.845 325.535 56.865 ;
        RECT 324.255 49.385 325.065 53.395 ;
        RECT 323.815 41.085 325.515 49.385 ;
        RECT 323.815 19.685 325.515 27.985 ;
        RECT 324.265 15.660 325.075 19.685 ;
        RECT 323.795 12.190 325.545 14.210 ;
        RECT 327.640 12.190 328.010 59.695 ;
        RECT 323.795 9.675 328.010 12.190 ;
        RECT 328.860 59.685 329.240 59.695 ;
        RECT 330.380 59.685 330.760 59.695 ;
        RECT 328.860 9.675 330.760 59.685 ;
        RECT 331.610 12.190 331.980 59.695 ;
        RECT 338.375 59.605 339.075 60.305 ;
        RECT 342.535 59.605 343.235 60.305 ;
        RECT 334.080 56.865 338.295 59.380 ;
        RECT 334.080 54.845 335.830 56.865 ;
        RECT 334.550 49.385 335.360 53.395 ;
        RECT 334.115 38.385 335.815 49.385 ;
        RECT 334.115 19.685 335.815 30.685 ;
        RECT 334.545 15.660 335.355 19.685 ;
        RECT 334.075 12.190 335.825 14.210 ;
        RECT 331.610 9.675 335.825 12.190 ;
        RECT 328.090 8.750 328.790 9.450 ;
        RECT 330.830 8.750 331.530 9.450 ;
        RECT 337.925 9.360 338.295 56.865 ;
        RECT 339.145 9.370 340.315 59.380 ;
        RECT 341.295 9.370 342.465 59.380 ;
        RECT 339.145 9.360 339.525 9.370 ;
        RECT 342.085 9.360 342.465 9.370 ;
        RECT 343.315 56.865 347.530 59.380 ;
        RECT 343.315 9.360 343.685 56.865 ;
        RECT 345.780 54.845 347.530 56.865 ;
        RECT 346.250 49.385 347.060 53.395 ;
        RECT 345.810 46.485 347.510 49.385 ;
        RECT 345.810 19.685 347.510 22.585 ;
        RECT 346.260 15.660 347.070 19.685 ;
        RECT 345.790 12.190 347.540 14.210 ;
        RECT 349.635 12.190 350.005 59.695 ;
        RECT 345.790 9.675 350.005 12.190 ;
        RECT 350.855 59.685 351.235 59.695 ;
        RECT 352.375 59.685 352.755 59.695 ;
        RECT 350.855 9.675 352.755 59.685 ;
        RECT 353.605 12.190 353.975 59.695 ;
        RECT 360.370 59.605 361.070 60.305 ;
        RECT 363.110 59.605 363.810 60.305 ;
        RECT 356.075 56.865 360.290 59.380 ;
        RECT 356.075 54.845 357.825 56.865 ;
        RECT 356.545 49.385 357.355 53.395 ;
        RECT 356.110 43.785 357.810 49.385 ;
        RECT 356.110 19.685 357.810 25.285 ;
        RECT 356.540 15.660 357.350 19.685 ;
        RECT 356.070 12.190 357.820 14.210 ;
        RECT 353.605 9.675 357.820 12.190 ;
        RECT 350.085 8.750 350.785 9.450 ;
        RECT 352.825 8.750 353.525 9.450 ;
        RECT 359.920 9.360 360.290 56.865 ;
        RECT 361.140 9.370 363.040 59.380 ;
        RECT 361.140 9.360 361.520 9.370 ;
        RECT 362.660 9.360 363.040 9.370 ;
        RECT 363.890 56.865 368.105 59.380 ;
        RECT 363.890 9.360 364.260 56.865 ;
        RECT 366.355 54.845 368.105 56.865 ;
        RECT 366.825 49.385 367.635 53.395 ;
        RECT 366.385 41.085 368.085 49.385 ;
        RECT 366.385 19.685 368.085 27.985 ;
        RECT 366.835 15.660 367.645 19.685 ;
        RECT 366.365 12.190 368.115 14.210 ;
        RECT 370.210 12.190 370.580 59.695 ;
        RECT 366.365 9.675 370.580 12.190 ;
        RECT 371.430 59.685 371.810 59.695 ;
        RECT 372.950 59.685 373.330 59.695 ;
        RECT 371.430 9.675 373.330 59.685 ;
        RECT 374.180 12.190 374.550 59.695 ;
        RECT 380.945 59.605 381.645 60.305 ;
        RECT 385.105 59.605 385.805 60.305 ;
        RECT 376.650 56.865 380.865 59.380 ;
        RECT 376.650 54.845 378.400 56.865 ;
        RECT 377.120 49.385 377.930 53.395 ;
        RECT 376.685 38.385 378.385 49.385 ;
        RECT 376.685 19.685 378.385 30.685 ;
        RECT 377.115 15.660 377.925 19.685 ;
        RECT 376.645 12.190 378.395 14.210 ;
        RECT 374.180 9.675 378.395 12.190 ;
        RECT 370.660 8.750 371.360 9.450 ;
        RECT 373.400 8.750 374.100 9.450 ;
        RECT 380.495 9.360 380.865 56.865 ;
        RECT 381.715 9.370 382.885 59.380 ;
        RECT 383.865 9.370 385.035 59.380 ;
        RECT 381.715 9.360 382.095 9.370 ;
        RECT 384.655 9.360 385.035 9.370 ;
        RECT 385.885 56.865 390.100 59.380 ;
        RECT 385.885 9.360 386.255 56.865 ;
        RECT 388.350 54.845 390.100 56.865 ;
        RECT 388.820 49.385 389.630 53.395 ;
        RECT 388.380 46.485 390.080 49.385 ;
        RECT 388.380 19.685 390.080 22.585 ;
        RECT 388.830 15.660 389.640 19.685 ;
        RECT 388.360 12.190 390.110 14.210 ;
        RECT 392.205 12.190 392.575 59.695 ;
        RECT 388.360 9.675 392.575 12.190 ;
        RECT 393.425 59.685 393.805 59.695 ;
        RECT 394.945 59.685 395.325 59.695 ;
        RECT 393.425 9.675 395.325 59.685 ;
        RECT 396.175 12.190 396.545 59.695 ;
        RECT 402.940 59.605 403.640 60.305 ;
        RECT 405.680 59.605 406.380 60.305 ;
        RECT 398.645 56.865 402.860 59.380 ;
        RECT 398.645 54.845 400.395 56.865 ;
        RECT 399.115 49.385 399.925 53.395 ;
        RECT 398.680 43.785 400.380 49.385 ;
        RECT 398.680 19.685 400.380 25.285 ;
        RECT 399.110 15.660 399.920 19.685 ;
        RECT 398.640 12.190 400.390 14.210 ;
        RECT 396.175 9.675 400.390 12.190 ;
        RECT 392.655 8.750 393.355 9.450 ;
        RECT 395.395 8.750 396.095 9.450 ;
        RECT 402.490 9.360 402.860 56.865 ;
        RECT 403.710 9.370 405.610 59.380 ;
        RECT 403.710 9.360 404.090 9.370 ;
        RECT 405.230 9.360 405.610 9.370 ;
        RECT 406.460 56.865 410.675 59.380 ;
        RECT 406.460 9.360 406.830 56.865 ;
        RECT 408.925 54.845 410.675 56.865 ;
        RECT 409.395 49.385 410.205 53.395 ;
        RECT 408.955 41.085 410.655 49.385 ;
        RECT 408.955 19.685 410.655 27.985 ;
        RECT 409.405 15.660 410.215 19.685 ;
        RECT 408.935 12.190 410.685 14.210 ;
        RECT 412.780 12.190 413.150 59.695 ;
        RECT 408.935 9.675 413.150 12.190 ;
        RECT 414.000 59.685 414.380 59.695 ;
        RECT 415.520 59.685 415.900 59.695 ;
        RECT 414.000 9.675 415.900 59.685 ;
        RECT 416.750 12.190 417.120 59.695 ;
        RECT 423.515 59.605 424.215 60.305 ;
        RECT 427.675 59.605 428.375 60.305 ;
        RECT 419.220 56.865 423.435 59.380 ;
        RECT 419.220 54.845 420.970 56.865 ;
        RECT 419.690 49.385 420.500 53.395 ;
        RECT 419.255 38.385 420.955 49.385 ;
        RECT 419.255 19.685 420.955 30.685 ;
        RECT 419.685 15.660 420.495 19.685 ;
        RECT 419.215 12.190 420.965 14.210 ;
        RECT 416.750 9.675 420.965 12.190 ;
        RECT 413.230 8.750 413.930 9.450 ;
        RECT 415.970 8.750 416.670 9.450 ;
        RECT 423.065 9.360 423.435 56.865 ;
        RECT 424.285 9.370 425.455 59.380 ;
        RECT 426.435 9.370 427.605 59.380 ;
        RECT 424.285 9.360 424.665 9.370 ;
        RECT 427.225 9.360 427.605 9.370 ;
        RECT 428.455 56.865 432.670 59.380 ;
        RECT 428.455 9.360 428.825 56.865 ;
        RECT 430.920 54.845 432.670 56.865 ;
        RECT 431.390 49.385 432.200 53.395 ;
        RECT 430.950 46.485 432.650 49.385 ;
        RECT 430.950 19.685 432.650 22.585 ;
        RECT 431.400 15.660 432.210 19.685 ;
        RECT 430.930 12.190 432.680 14.210 ;
        RECT 434.775 12.190 435.145 59.695 ;
        RECT 430.930 9.675 435.145 12.190 ;
        RECT 435.995 59.685 436.375 59.695 ;
        RECT 437.515 59.685 437.895 59.695 ;
        RECT 435.995 9.675 437.895 59.685 ;
        RECT 438.745 12.190 439.115 59.695 ;
        RECT 445.510 59.605 446.210 60.305 ;
        RECT 448.250 59.605 448.950 60.305 ;
        RECT 441.215 56.865 445.430 59.380 ;
        RECT 441.215 54.845 442.965 56.865 ;
        RECT 441.685 49.385 442.495 53.395 ;
        RECT 441.250 43.785 442.950 49.385 ;
        RECT 441.250 19.685 442.950 25.285 ;
        RECT 441.680 15.660 442.490 19.685 ;
        RECT 441.210 12.190 442.960 14.210 ;
        RECT 438.745 9.675 442.960 12.190 ;
        RECT 435.225 8.750 435.925 9.450 ;
        RECT 437.965 8.750 438.665 9.450 ;
        RECT 445.060 9.360 445.430 56.865 ;
        RECT 446.280 9.370 448.180 59.380 ;
        RECT 446.280 9.360 446.660 9.370 ;
        RECT 447.800 9.360 448.180 9.370 ;
        RECT 449.030 56.865 453.245 59.380 ;
        RECT 449.030 9.360 449.400 56.865 ;
        RECT 451.495 54.845 453.245 56.865 ;
        RECT 451.965 49.385 452.775 53.395 ;
        RECT 451.525 41.085 453.225 49.385 ;
        RECT 451.525 19.685 453.225 27.985 ;
        RECT 451.975 15.660 452.785 19.685 ;
        RECT 451.505 12.190 453.255 14.210 ;
        RECT 455.350 12.190 455.720 59.695 ;
        RECT 451.505 9.675 455.720 12.190 ;
        RECT 456.570 59.685 456.950 59.695 ;
        RECT 458.090 59.685 458.470 59.695 ;
        RECT 456.570 9.675 458.470 59.685 ;
        RECT 459.320 12.190 459.690 59.695 ;
        RECT 466.085 59.605 466.785 60.305 ;
        RECT 470.245 59.605 470.945 60.305 ;
        RECT 461.790 56.865 466.005 59.380 ;
        RECT 461.790 54.845 463.540 56.865 ;
        RECT 462.260 49.385 463.070 53.395 ;
        RECT 461.825 38.385 463.525 49.385 ;
        RECT 461.825 19.685 463.525 30.685 ;
        RECT 462.255 15.660 463.065 19.685 ;
        RECT 461.785 12.190 463.535 14.210 ;
        RECT 459.320 9.675 463.535 12.190 ;
        RECT 455.800 8.750 456.500 9.450 ;
        RECT 458.540 8.750 459.240 9.450 ;
        RECT 465.635 9.360 466.005 56.865 ;
        RECT 466.855 9.370 468.025 59.380 ;
        RECT 469.005 9.370 470.175 59.380 ;
        RECT 466.855 9.360 467.235 9.370 ;
        RECT 469.795 9.360 470.175 9.370 ;
        RECT 471.025 56.865 475.240 59.380 ;
        RECT 471.025 9.360 471.395 56.865 ;
        RECT 473.490 54.845 475.240 56.865 ;
        RECT 473.960 49.385 474.770 53.395 ;
        RECT 473.520 46.485 475.220 49.385 ;
        RECT 473.520 19.685 475.220 22.585 ;
        RECT 473.970 15.660 474.780 19.685 ;
        RECT 473.500 12.190 475.250 14.210 ;
        RECT 477.345 12.190 477.715 59.695 ;
        RECT 473.500 9.675 477.715 12.190 ;
        RECT 478.565 59.685 478.945 59.695 ;
        RECT 480.085 59.685 480.465 59.695 ;
        RECT 478.565 9.675 480.465 59.685 ;
        RECT 481.315 12.190 481.685 59.695 ;
        RECT 488.080 59.605 488.780 60.305 ;
        RECT 490.820 59.605 491.520 60.305 ;
        RECT 483.785 56.865 488.000 59.380 ;
        RECT 483.785 54.845 485.535 56.865 ;
        RECT 484.255 49.385 485.065 53.395 ;
        RECT 483.820 43.785 485.520 49.385 ;
        RECT 483.820 19.685 485.520 25.285 ;
        RECT 484.250 15.660 485.060 19.685 ;
        RECT 483.780 12.190 485.530 14.210 ;
        RECT 481.315 9.675 485.530 12.190 ;
        RECT 477.795 8.750 478.495 9.450 ;
        RECT 480.535 8.750 481.235 9.450 ;
        RECT 487.630 9.360 488.000 56.865 ;
        RECT 488.850 9.370 490.750 59.380 ;
        RECT 488.850 9.360 489.230 9.370 ;
        RECT 490.370 9.360 490.750 9.370 ;
        RECT 491.600 56.865 495.815 59.380 ;
        RECT 491.600 9.360 491.970 56.865 ;
        RECT 494.065 54.845 495.815 56.865 ;
        RECT 494.535 49.385 495.345 53.395 ;
        RECT 494.095 41.085 495.795 49.385 ;
        RECT 494.095 19.685 495.795 27.985 ;
        RECT 494.545 15.660 495.355 19.685 ;
        RECT 494.075 12.190 495.825 14.210 ;
        RECT 497.920 12.190 498.290 59.695 ;
        RECT 494.075 9.675 498.290 12.190 ;
        RECT 499.140 59.685 499.520 59.695 ;
        RECT 500.660 59.685 501.040 59.695 ;
        RECT 499.140 9.675 501.040 59.685 ;
        RECT 501.890 12.190 502.260 59.695 ;
        RECT 508.655 59.605 509.355 60.305 ;
        RECT 512.815 59.605 513.515 60.305 ;
        RECT 504.360 56.865 508.575 59.380 ;
        RECT 504.360 54.845 506.110 56.865 ;
        RECT 504.830 49.385 505.640 53.395 ;
        RECT 504.395 38.385 506.095 49.385 ;
        RECT 504.395 19.685 506.095 30.685 ;
        RECT 504.825 15.660 505.635 19.685 ;
        RECT 504.355 12.190 506.105 14.210 ;
        RECT 501.890 9.675 506.105 12.190 ;
        RECT 498.370 8.750 499.070 9.450 ;
        RECT 501.110 8.750 501.810 9.450 ;
        RECT 508.205 9.360 508.575 56.865 ;
        RECT 509.425 9.370 510.595 59.380 ;
        RECT 511.575 9.370 512.745 59.380 ;
        RECT 509.425 9.360 509.805 9.370 ;
        RECT 512.365 9.360 512.745 9.370 ;
        RECT 513.595 56.865 517.810 59.380 ;
        RECT 513.595 9.360 513.965 56.865 ;
        RECT 516.060 54.845 517.810 56.865 ;
        RECT 516.530 49.385 517.340 53.395 ;
        RECT 516.090 46.485 517.790 49.385 ;
        RECT 516.090 19.685 517.790 22.585 ;
        RECT 516.540 15.660 517.350 19.685 ;
        RECT 516.070 12.190 517.820 14.210 ;
        RECT 519.915 12.190 520.285 59.695 ;
        RECT 516.070 9.675 520.285 12.190 ;
        RECT 521.135 59.685 521.515 59.695 ;
        RECT 522.655 59.685 523.035 59.695 ;
        RECT 521.135 9.675 523.035 59.685 ;
        RECT 523.885 12.190 524.255 59.695 ;
        RECT 530.650 59.605 531.350 60.305 ;
        RECT 533.390 59.605 534.090 60.305 ;
        RECT 526.355 56.865 530.570 59.380 ;
        RECT 526.355 54.845 528.105 56.865 ;
        RECT 526.825 49.385 527.635 53.395 ;
        RECT 526.390 43.785 528.090 49.385 ;
        RECT 526.390 19.685 528.090 25.285 ;
        RECT 526.820 15.660 527.630 19.685 ;
        RECT 526.350 12.190 528.100 14.210 ;
        RECT 523.885 9.675 528.100 12.190 ;
        RECT 520.365 8.750 521.065 9.450 ;
        RECT 523.105 8.750 523.805 9.450 ;
        RECT 530.200 9.360 530.570 56.865 ;
        RECT 531.420 9.370 533.320 59.380 ;
        RECT 531.420 9.360 531.800 9.370 ;
        RECT 532.940 9.360 533.320 9.370 ;
        RECT 534.170 56.865 538.385 59.380 ;
        RECT 534.170 9.360 534.540 56.865 ;
        RECT 536.635 54.845 538.385 56.865 ;
        RECT 537.105 49.385 537.915 53.395 ;
        RECT 536.665 41.085 538.365 49.385 ;
        RECT 536.665 19.685 538.365 27.985 ;
        RECT 537.115 15.660 537.925 19.685 ;
        RECT 536.645 12.190 538.395 14.210 ;
        RECT 540.490 12.190 540.860 59.695 ;
        RECT 536.645 9.675 540.860 12.190 ;
        RECT 541.710 59.685 542.090 59.695 ;
        RECT 543.230 59.685 543.610 59.695 ;
        RECT 541.710 9.675 543.610 59.685 ;
        RECT 544.460 12.190 544.830 59.695 ;
        RECT 551.225 59.605 551.925 60.305 ;
        RECT 555.385 59.605 556.085 60.305 ;
        RECT 546.930 56.865 551.145 59.380 ;
        RECT 546.930 54.845 548.680 56.865 ;
        RECT 547.400 49.385 548.210 53.395 ;
        RECT 546.965 38.385 548.665 49.385 ;
        RECT 546.965 19.685 548.665 30.685 ;
        RECT 547.395 15.660 548.205 19.685 ;
        RECT 546.925 12.190 548.675 14.210 ;
        RECT 544.460 9.675 548.675 12.190 ;
        RECT 540.940 8.750 541.640 9.450 ;
        RECT 543.680 8.750 544.380 9.450 ;
        RECT 550.775 9.360 551.145 56.865 ;
        RECT 551.995 9.370 553.165 59.380 ;
        RECT 554.145 9.370 555.315 59.380 ;
        RECT 551.995 9.360 552.375 9.370 ;
        RECT 554.935 9.360 555.315 9.370 ;
        RECT 556.165 56.865 560.380 59.380 ;
        RECT 556.165 9.360 556.535 56.865 ;
        RECT 558.630 54.845 560.380 56.865 ;
        RECT 559.100 49.385 559.910 53.395 ;
        RECT 558.660 46.485 560.360 49.385 ;
        RECT 558.660 19.685 560.360 22.585 ;
        RECT 559.110 15.660 559.920 19.685 ;
        RECT 558.640 12.190 560.390 14.210 ;
        RECT 562.485 12.190 562.855 59.695 ;
        RECT 558.640 9.675 562.855 12.190 ;
        RECT 563.705 59.685 564.085 59.695 ;
        RECT 565.225 59.685 565.605 59.695 ;
        RECT 563.705 9.675 565.605 59.685 ;
        RECT 566.455 12.190 566.825 59.695 ;
        RECT 573.220 59.605 573.920 60.305 ;
        RECT 575.960 59.605 576.660 60.305 ;
        RECT 568.925 56.865 573.140 59.380 ;
        RECT 568.925 54.845 570.675 56.865 ;
        RECT 569.395 49.385 570.205 53.395 ;
        RECT 568.960 43.785 570.660 49.385 ;
        RECT 568.960 19.685 570.660 25.285 ;
        RECT 569.390 15.660 570.200 19.685 ;
        RECT 568.920 12.190 570.670 14.210 ;
        RECT 566.455 9.675 570.670 12.190 ;
        RECT 562.935 8.750 563.635 9.450 ;
        RECT 565.675 8.750 566.375 9.450 ;
        RECT 572.770 9.360 573.140 56.865 ;
        RECT 573.990 9.370 575.890 59.380 ;
        RECT 573.990 9.360 574.370 9.370 ;
        RECT 575.510 9.360 575.890 9.370 ;
        RECT 576.740 56.865 580.955 59.380 ;
        RECT 576.740 9.360 577.110 56.865 ;
        RECT 579.205 54.845 580.955 56.865 ;
        RECT 579.675 49.385 580.485 53.395 ;
        RECT 579.235 41.085 580.935 49.385 ;
        RECT 579.235 19.685 580.935 27.985 ;
        RECT 579.685 15.660 580.495 19.685 ;
        RECT 579.215 12.190 580.965 14.210 ;
        RECT 583.060 12.190 583.430 59.695 ;
        RECT 579.215 9.675 583.430 12.190 ;
        RECT 584.280 59.685 584.660 59.695 ;
        RECT 585.800 59.685 586.180 59.695 ;
        RECT 584.280 9.675 586.180 59.685 ;
        RECT 587.030 12.190 587.400 59.695 ;
        RECT 593.795 59.605 594.495 60.305 ;
        RECT 597.955 59.605 598.655 60.305 ;
        RECT 589.500 56.865 593.715 59.380 ;
        RECT 589.500 54.845 591.250 56.865 ;
        RECT 589.970 49.385 590.780 53.395 ;
        RECT 589.535 38.385 591.235 49.385 ;
        RECT 589.535 19.685 591.235 30.685 ;
        RECT 589.965 15.660 590.775 19.685 ;
        RECT 589.495 12.190 591.245 14.210 ;
        RECT 587.030 9.675 591.245 12.190 ;
        RECT 583.510 8.750 584.210 9.450 ;
        RECT 586.250 8.750 586.950 9.450 ;
        RECT 593.345 9.360 593.715 56.865 ;
        RECT 594.565 9.370 595.735 59.380 ;
        RECT 596.715 9.370 597.885 59.380 ;
        RECT 594.565 9.360 594.945 9.370 ;
        RECT 597.505 9.360 597.885 9.370 ;
        RECT 598.735 56.865 602.950 59.380 ;
        RECT 598.735 9.360 599.105 56.865 ;
        RECT 601.200 54.845 602.950 56.865 ;
        RECT 601.670 49.385 602.480 53.395 ;
        RECT 601.230 46.485 602.930 49.385 ;
        RECT 601.230 19.685 602.930 22.585 ;
        RECT 601.680 15.660 602.490 19.685 ;
        RECT 601.210 12.190 602.960 14.210 ;
        RECT 605.055 12.190 605.425 59.695 ;
        RECT 601.210 9.675 605.425 12.190 ;
        RECT 606.275 59.685 606.655 59.695 ;
        RECT 607.795 59.685 608.175 59.695 ;
        RECT 606.275 9.675 608.175 59.685 ;
        RECT 609.025 12.190 609.395 59.695 ;
        RECT 615.790 59.605 616.490 60.305 ;
        RECT 618.530 59.605 619.230 60.305 ;
        RECT 611.495 56.865 615.710 59.380 ;
        RECT 611.495 54.845 613.245 56.865 ;
        RECT 611.965 49.385 612.775 53.395 ;
        RECT 611.530 43.785 613.230 49.385 ;
        RECT 611.530 19.685 613.230 25.285 ;
        RECT 611.960 15.660 612.770 19.685 ;
        RECT 611.490 12.190 613.240 14.210 ;
        RECT 609.025 9.675 613.240 12.190 ;
        RECT 605.505 8.750 606.205 9.450 ;
        RECT 608.245 8.750 608.945 9.450 ;
        RECT 615.340 9.360 615.710 56.865 ;
        RECT 616.560 9.370 618.460 59.380 ;
        RECT 616.560 9.360 616.940 9.370 ;
        RECT 618.080 9.360 618.460 9.370 ;
        RECT 619.310 56.865 623.525 59.380 ;
        RECT 619.310 9.360 619.680 56.865 ;
        RECT 621.775 54.845 623.525 56.865 ;
        RECT 622.245 49.385 623.055 53.395 ;
        RECT 621.805 41.085 623.505 49.385 ;
        RECT 621.805 19.685 623.505 27.985 ;
        RECT 622.255 15.660 623.065 19.685 ;
        RECT 621.785 12.190 623.535 14.210 ;
        RECT 625.630 12.190 626.000 59.695 ;
        RECT 621.785 9.675 626.000 12.190 ;
        RECT 626.850 59.685 627.230 59.695 ;
        RECT 628.370 59.685 628.750 59.695 ;
        RECT 626.850 9.675 628.750 59.685 ;
        RECT 629.600 12.190 629.970 59.695 ;
        RECT 636.365 59.605 637.065 60.305 ;
        RECT 640.525 59.605 641.225 60.305 ;
        RECT 632.070 56.865 636.285 59.380 ;
        RECT 632.070 54.845 633.820 56.865 ;
        RECT 632.540 49.385 633.350 53.395 ;
        RECT 632.105 38.385 633.805 49.385 ;
        RECT 632.105 19.685 633.805 30.685 ;
        RECT 632.535 15.660 633.345 19.685 ;
        RECT 632.065 12.190 633.815 14.210 ;
        RECT 629.600 9.675 633.815 12.190 ;
        RECT 626.080 8.750 626.780 9.450 ;
        RECT 628.820 8.750 629.520 9.450 ;
        RECT 635.915 9.360 636.285 56.865 ;
        RECT 637.135 9.370 638.305 59.380 ;
        RECT 639.285 9.370 640.455 59.380 ;
        RECT 637.135 9.360 637.515 9.370 ;
        RECT 640.075 9.360 640.455 9.370 ;
        RECT 641.305 56.865 645.520 59.380 ;
        RECT 641.305 9.360 641.675 56.865 ;
        RECT 643.770 54.845 645.520 56.865 ;
        RECT 644.240 49.385 645.050 53.395 ;
        RECT 643.800 46.485 645.500 49.385 ;
        RECT 643.800 19.685 645.500 22.585 ;
        RECT 644.250 15.660 645.060 19.685 ;
        RECT 643.780 12.190 645.530 14.210 ;
        RECT 647.625 12.190 647.995 59.695 ;
        RECT 643.780 9.675 647.995 12.190 ;
        RECT 648.845 59.685 649.225 59.695 ;
        RECT 650.365 59.685 650.745 59.695 ;
        RECT 648.845 9.675 650.745 59.685 ;
        RECT 651.595 12.190 651.965 59.695 ;
        RECT 658.360 59.605 659.060 60.305 ;
        RECT 661.100 59.605 661.800 60.305 ;
        RECT 654.065 56.865 658.280 59.380 ;
        RECT 654.065 54.845 655.815 56.865 ;
        RECT 654.535 49.385 655.345 53.395 ;
        RECT 654.100 43.785 655.800 49.385 ;
        RECT 654.100 19.685 655.800 25.285 ;
        RECT 654.530 15.660 655.340 19.685 ;
        RECT 654.060 12.190 655.810 14.210 ;
        RECT 651.595 9.675 655.810 12.190 ;
        RECT 648.075 8.750 648.775 9.450 ;
        RECT 650.815 8.750 651.515 9.450 ;
        RECT 657.910 9.360 658.280 56.865 ;
        RECT 659.130 9.370 661.030 59.380 ;
        RECT 659.130 9.360 659.510 9.370 ;
        RECT 660.650 9.360 661.030 9.370 ;
        RECT 661.880 56.865 666.095 59.380 ;
        RECT 661.880 9.360 662.250 56.865 ;
        RECT 664.345 54.845 666.095 56.865 ;
        RECT 664.815 49.385 665.625 53.395 ;
        RECT 664.375 41.085 666.075 49.385 ;
        RECT 664.375 19.685 666.075 27.985 ;
        RECT 664.825 15.660 665.635 19.685 ;
        RECT 664.355 12.190 666.105 14.210 ;
        RECT 668.200 12.190 668.570 59.695 ;
        RECT 664.355 9.675 668.570 12.190 ;
        RECT 669.420 59.685 669.800 59.695 ;
        RECT 670.940 59.685 671.320 59.695 ;
        RECT 669.420 9.675 671.320 59.685 ;
        RECT 672.170 12.190 672.540 59.695 ;
        RECT 678.935 59.605 679.635 60.305 ;
        RECT 674.640 56.865 678.855 59.380 ;
        RECT 674.640 54.845 676.390 56.865 ;
        RECT 675.110 49.385 675.920 53.395 ;
        RECT 674.675 38.385 676.375 49.385 ;
        RECT 674.675 19.685 676.375 30.685 ;
        RECT 675.105 15.660 675.915 19.685 ;
        RECT 674.635 12.190 676.385 14.210 ;
        RECT 672.170 9.675 676.385 12.190 ;
        RECT 668.650 8.750 669.350 9.450 ;
        RECT 671.390 8.750 672.090 9.450 ;
        RECT 678.485 9.360 678.855 56.865 ;
        RECT 679.705 9.370 680.875 59.380 ;
        RECT 679.705 9.360 680.085 9.370 ;
        RECT 682.280 9.185 682.720 59.185 ;
        RECT 682.310 8.875 682.690 9.185 ;
        RECT 683.070 9.175 683.450 59.195 ;
        RECT 684.100 55.495 684.470 59.195 ;
        RECT 684.095 55.115 684.475 55.495 ;
        RECT 684.100 54.835 684.470 55.115 ;
        RECT 684.095 54.455 684.475 54.835 ;
        RECT 684.100 54.175 684.470 54.455 ;
        RECT 684.095 53.795 684.475 54.175 ;
        RECT 684.100 53.515 684.470 53.795 ;
        RECT 684.095 53.135 684.475 53.515 ;
        RECT 684.100 52.855 684.470 53.135 ;
        RECT 684.095 52.475 684.475 52.855 ;
        RECT 684.100 52.195 684.470 52.475 ;
        RECT 684.095 51.815 684.475 52.195 ;
        RECT 684.100 51.535 684.470 51.815 ;
        RECT 684.095 51.155 684.475 51.535 ;
        RECT 684.100 50.875 684.470 51.155 ;
        RECT 684.095 50.495 684.475 50.875 ;
        RECT 684.100 18.495 684.470 50.495 ;
        RECT 684.095 18.115 684.475 18.495 ;
        RECT 684.100 17.835 684.470 18.115 ;
        RECT 684.095 17.455 684.475 17.835 ;
        RECT 684.100 17.175 684.470 17.455 ;
        RECT 684.095 16.795 684.475 17.175 ;
        RECT 684.100 16.515 684.470 16.795 ;
        RECT 684.095 16.135 684.475 16.515 ;
        RECT 684.100 15.855 684.470 16.135 ;
        RECT 684.095 15.475 684.475 15.855 ;
        RECT 684.100 15.195 684.470 15.475 ;
        RECT 684.095 14.815 684.475 15.195 ;
        RECT 684.100 14.535 684.470 14.815 ;
        RECT 684.095 14.155 684.475 14.535 ;
        RECT 684.100 13.875 684.470 14.155 ;
        RECT 684.095 13.495 684.475 13.875 ;
        RECT 684.100 13.215 684.470 13.495 ;
        RECT 684.095 12.835 684.475 13.215 ;
        RECT 684.100 12.555 684.470 12.835 ;
        RECT 684.095 12.175 684.475 12.555 ;
        RECT 684.100 11.895 684.470 12.175 ;
        RECT 684.095 11.515 684.475 11.895 ;
        RECT 684.100 11.235 684.470 11.515 ;
        RECT 684.095 10.855 684.475 11.235 ;
        RECT 684.100 10.575 684.470 10.855 ;
        RECT 684.095 10.195 684.475 10.575 ;
        RECT 684.100 9.915 684.470 10.195 ;
        RECT 684.095 9.535 684.475 9.915 ;
        RECT 684.100 9.255 684.470 9.535 ;
        RECT 684.095 8.875 684.475 9.255 ;
        RECT 686.920 9.185 687.360 59.185 ;
        RECT 686.950 8.875 687.330 9.185 ;
        RECT 687.710 9.175 688.090 59.195 ;
        RECT 688.740 55.495 689.110 59.195 ;
        RECT 688.735 55.115 689.115 55.495 ;
        RECT 688.740 54.835 689.110 55.115 ;
        RECT 688.735 54.455 689.115 54.835 ;
        RECT 688.740 54.175 689.110 54.455 ;
        RECT 688.735 53.795 689.115 54.175 ;
        RECT 688.740 53.515 689.110 53.795 ;
        RECT 688.735 53.135 689.115 53.515 ;
        RECT 688.740 52.855 689.110 53.135 ;
        RECT 688.735 52.475 689.115 52.855 ;
        RECT 688.740 52.195 689.110 52.475 ;
        RECT 688.735 51.815 689.115 52.195 ;
        RECT 688.740 51.535 689.110 51.815 ;
        RECT 688.735 51.155 689.115 51.535 ;
        RECT 688.740 50.875 689.110 51.155 ;
        RECT 688.735 50.495 689.115 50.875 ;
        RECT 688.740 18.495 689.110 50.495 ;
        RECT 688.735 18.115 689.115 18.495 ;
        RECT 688.740 17.835 689.110 18.115 ;
        RECT 688.735 17.455 689.115 17.835 ;
        RECT 688.740 17.175 689.110 17.455 ;
        RECT 688.735 16.795 689.115 17.175 ;
        RECT 688.740 16.515 689.110 16.795 ;
        RECT 688.735 16.135 689.115 16.515 ;
        RECT 688.740 15.855 689.110 16.135 ;
        RECT 688.735 15.475 689.115 15.855 ;
        RECT 688.740 15.195 689.110 15.475 ;
        RECT 688.735 14.815 689.115 15.195 ;
        RECT 688.740 14.535 689.110 14.815 ;
        RECT 688.735 14.155 689.115 14.535 ;
        RECT 688.740 13.875 689.110 14.155 ;
        RECT 688.735 13.495 689.115 13.875 ;
        RECT 688.740 13.215 689.110 13.495 ;
        RECT 688.735 12.835 689.115 13.215 ;
        RECT 688.740 12.555 689.110 12.835 ;
        RECT 688.735 12.175 689.115 12.555 ;
        RECT 688.740 11.895 689.110 12.175 ;
        RECT 688.735 11.515 689.115 11.895 ;
        RECT 688.740 11.235 689.110 11.515 ;
        RECT 688.735 10.855 689.115 11.235 ;
        RECT 688.740 10.575 689.110 10.855 ;
        RECT 688.735 10.195 689.115 10.575 ;
        RECT 688.740 9.915 689.110 10.195 ;
        RECT 688.735 9.535 689.115 9.915 ;
        RECT 688.740 9.255 689.110 9.535 ;
        RECT 688.735 8.875 689.115 9.255 ;
        RECT 691.560 9.185 692.000 59.185 ;
        RECT 691.590 8.875 691.970 9.185 ;
        RECT 692.350 9.175 692.730 59.195 ;
        RECT 693.380 55.495 693.750 59.195 ;
        RECT 693.375 55.115 693.755 55.495 ;
        RECT 693.380 54.835 693.750 55.115 ;
        RECT 693.375 54.455 693.755 54.835 ;
        RECT 693.380 54.175 693.750 54.455 ;
        RECT 693.375 53.795 693.755 54.175 ;
        RECT 693.380 53.515 693.750 53.795 ;
        RECT 693.375 53.135 693.755 53.515 ;
        RECT 693.380 52.855 693.750 53.135 ;
        RECT 693.375 52.475 693.755 52.855 ;
        RECT 693.380 52.195 693.750 52.475 ;
        RECT 693.375 51.815 693.755 52.195 ;
        RECT 693.380 51.535 693.750 51.815 ;
        RECT 693.375 51.155 693.755 51.535 ;
        RECT 693.380 50.875 693.750 51.155 ;
        RECT 693.375 50.495 693.755 50.875 ;
        RECT 693.380 18.495 693.750 50.495 ;
        RECT 693.375 18.115 693.755 18.495 ;
        RECT 693.380 17.835 693.750 18.115 ;
        RECT 693.375 17.455 693.755 17.835 ;
        RECT 693.380 17.175 693.750 17.455 ;
        RECT 693.375 16.795 693.755 17.175 ;
        RECT 693.380 16.515 693.750 16.795 ;
        RECT 693.375 16.135 693.755 16.515 ;
        RECT 693.380 15.855 693.750 16.135 ;
        RECT 693.375 15.475 693.755 15.855 ;
        RECT 693.380 15.195 693.750 15.475 ;
        RECT 693.375 14.815 693.755 15.195 ;
        RECT 693.380 14.535 693.750 14.815 ;
        RECT 693.375 14.155 693.755 14.535 ;
        RECT 693.380 13.875 693.750 14.155 ;
        RECT 693.375 13.495 693.755 13.875 ;
        RECT 693.380 13.215 693.750 13.495 ;
        RECT 693.375 12.835 693.755 13.215 ;
        RECT 693.380 12.555 693.750 12.835 ;
        RECT 693.375 12.175 693.755 12.555 ;
        RECT 693.380 11.895 693.750 12.175 ;
        RECT 693.375 11.515 693.755 11.895 ;
        RECT 693.380 11.235 693.750 11.515 ;
        RECT 693.375 10.855 693.755 11.235 ;
        RECT 693.380 10.575 693.750 10.855 ;
        RECT 693.375 10.195 693.755 10.575 ;
        RECT 693.380 9.915 693.750 10.195 ;
        RECT 693.375 9.535 693.755 9.915 ;
        RECT 693.380 9.255 693.750 9.535 ;
        RECT 693.375 8.875 693.755 9.255 ;
        RECT 696.200 9.185 696.640 59.185 ;
        RECT 696.230 8.875 696.610 9.185 ;
        RECT 696.990 9.175 697.370 59.195 ;
        RECT 698.020 55.495 698.390 59.195 ;
        RECT 698.015 55.115 698.395 55.495 ;
        RECT 698.020 54.835 698.390 55.115 ;
        RECT 698.015 54.455 698.395 54.835 ;
        RECT 698.020 54.175 698.390 54.455 ;
        RECT 698.015 53.795 698.395 54.175 ;
        RECT 698.020 53.515 698.390 53.795 ;
        RECT 698.015 53.135 698.395 53.515 ;
        RECT 698.020 52.855 698.390 53.135 ;
        RECT 698.015 52.475 698.395 52.855 ;
        RECT 698.020 52.195 698.390 52.475 ;
        RECT 698.015 51.815 698.395 52.195 ;
        RECT 698.020 51.535 698.390 51.815 ;
        RECT 698.015 51.155 698.395 51.535 ;
        RECT 698.020 50.875 698.390 51.155 ;
        RECT 698.015 50.495 698.395 50.875 ;
        RECT 698.020 18.495 698.390 50.495 ;
        RECT 698.015 18.115 698.395 18.495 ;
        RECT 698.020 17.835 698.390 18.115 ;
        RECT 698.015 17.455 698.395 17.835 ;
        RECT 698.020 17.175 698.390 17.455 ;
        RECT 698.015 16.795 698.395 17.175 ;
        RECT 698.020 16.515 698.390 16.795 ;
        RECT 698.015 16.135 698.395 16.515 ;
        RECT 698.020 15.855 698.390 16.135 ;
        RECT 698.015 15.475 698.395 15.855 ;
        RECT 698.020 15.195 698.390 15.475 ;
        RECT 698.015 14.815 698.395 15.195 ;
        RECT 698.020 14.535 698.390 14.815 ;
        RECT 698.015 14.155 698.395 14.535 ;
        RECT 698.020 13.875 698.390 14.155 ;
        RECT 698.015 13.495 698.395 13.875 ;
        RECT 698.020 13.215 698.390 13.495 ;
        RECT 698.015 12.835 698.395 13.215 ;
        RECT 698.020 12.555 698.390 12.835 ;
        RECT 698.015 12.175 698.395 12.555 ;
        RECT 698.020 11.895 698.390 12.175 ;
        RECT 698.015 11.515 698.395 11.895 ;
        RECT 698.020 11.235 698.390 11.515 ;
        RECT 698.015 10.855 698.395 11.235 ;
        RECT 698.020 10.575 698.390 10.855 ;
        RECT 698.015 10.195 698.395 10.575 ;
        RECT 698.020 9.915 698.390 10.195 ;
        RECT 698.015 9.535 698.395 9.915 ;
        RECT 698.020 9.255 698.390 9.535 ;
        RECT 698.015 8.875 698.395 9.255 ;
        RECT 700.840 9.185 701.280 59.185 ;
        RECT 700.870 8.875 701.250 9.185 ;
        RECT 701.630 9.175 702.010 59.195 ;
        RECT 702.660 55.495 703.030 59.195 ;
        RECT 702.655 55.115 703.035 55.495 ;
        RECT 702.660 54.835 703.030 55.115 ;
        RECT 702.655 54.455 703.035 54.835 ;
        RECT 702.660 54.175 703.030 54.455 ;
        RECT 702.655 53.795 703.035 54.175 ;
        RECT 702.660 53.515 703.030 53.795 ;
        RECT 702.655 53.135 703.035 53.515 ;
        RECT 702.660 52.855 703.030 53.135 ;
        RECT 702.655 52.475 703.035 52.855 ;
        RECT 702.660 52.195 703.030 52.475 ;
        RECT 702.655 51.815 703.035 52.195 ;
        RECT 702.660 51.535 703.030 51.815 ;
        RECT 702.655 51.155 703.035 51.535 ;
        RECT 702.660 50.875 703.030 51.155 ;
        RECT 702.655 50.495 703.035 50.875 ;
        RECT 702.660 18.495 703.030 50.495 ;
        RECT 702.655 18.115 703.035 18.495 ;
        RECT 702.660 17.835 703.030 18.115 ;
        RECT 702.655 17.455 703.035 17.835 ;
        RECT 702.660 17.175 703.030 17.455 ;
        RECT 702.655 16.795 703.035 17.175 ;
        RECT 702.660 16.515 703.030 16.795 ;
        RECT 702.655 16.135 703.035 16.515 ;
        RECT 702.660 15.855 703.030 16.135 ;
        RECT 702.655 15.475 703.035 15.855 ;
        RECT 702.660 15.195 703.030 15.475 ;
        RECT 702.655 14.815 703.035 15.195 ;
        RECT 702.660 14.535 703.030 14.815 ;
        RECT 702.655 14.155 703.035 14.535 ;
        RECT 702.660 13.875 703.030 14.155 ;
        RECT 702.655 13.495 703.035 13.875 ;
        RECT 702.660 13.215 703.030 13.495 ;
        RECT 702.655 12.835 703.035 13.215 ;
        RECT 702.660 12.555 703.030 12.835 ;
        RECT 702.655 12.175 703.035 12.555 ;
        RECT 702.660 11.895 703.030 12.175 ;
        RECT 702.655 11.515 703.035 11.895 ;
        RECT 702.660 11.235 703.030 11.515 ;
        RECT 702.655 10.855 703.035 11.235 ;
        RECT 702.660 10.575 703.030 10.855 ;
        RECT 702.655 10.195 703.035 10.575 ;
        RECT 702.660 9.915 703.030 10.195 ;
        RECT 702.655 9.535 703.035 9.915 ;
        RECT 702.660 9.255 703.030 9.535 ;
        RECT 702.655 8.875 703.035 9.255 ;
        RECT 705.480 9.185 705.920 59.185 ;
        RECT 705.510 8.875 705.890 9.185 ;
        RECT 706.270 9.175 706.650 59.195 ;
        RECT 707.300 55.495 707.670 59.195 ;
        RECT 707.295 55.115 707.675 55.495 ;
        RECT 707.300 54.835 707.670 55.115 ;
        RECT 707.295 54.455 707.675 54.835 ;
        RECT 707.300 54.175 707.670 54.455 ;
        RECT 707.295 53.795 707.675 54.175 ;
        RECT 707.300 53.515 707.670 53.795 ;
        RECT 707.295 53.135 707.675 53.515 ;
        RECT 707.300 52.855 707.670 53.135 ;
        RECT 707.295 52.475 707.675 52.855 ;
        RECT 707.300 52.195 707.670 52.475 ;
        RECT 707.295 51.815 707.675 52.195 ;
        RECT 707.300 51.535 707.670 51.815 ;
        RECT 707.295 51.155 707.675 51.535 ;
        RECT 707.300 50.875 707.670 51.155 ;
        RECT 707.295 50.495 707.675 50.875 ;
        RECT 707.300 18.495 707.670 50.495 ;
        RECT 707.295 18.115 707.675 18.495 ;
        RECT 707.300 17.835 707.670 18.115 ;
        RECT 707.295 17.455 707.675 17.835 ;
        RECT 707.300 17.175 707.670 17.455 ;
        RECT 707.295 16.795 707.675 17.175 ;
        RECT 707.300 16.515 707.670 16.795 ;
        RECT 707.295 16.135 707.675 16.515 ;
        RECT 707.300 15.855 707.670 16.135 ;
        RECT 707.295 15.475 707.675 15.855 ;
        RECT 707.300 15.195 707.670 15.475 ;
        RECT 707.295 14.815 707.675 15.195 ;
        RECT 707.300 14.535 707.670 14.815 ;
        RECT 707.295 14.155 707.675 14.535 ;
        RECT 707.300 13.875 707.670 14.155 ;
        RECT 707.295 13.495 707.675 13.875 ;
        RECT 707.300 13.215 707.670 13.495 ;
        RECT 707.295 12.835 707.675 13.215 ;
        RECT 707.300 12.555 707.670 12.835 ;
        RECT 707.295 12.175 707.675 12.555 ;
        RECT 707.300 11.895 707.670 12.175 ;
        RECT 707.295 11.515 707.675 11.895 ;
        RECT 707.300 11.235 707.670 11.515 ;
        RECT 707.295 10.855 707.675 11.235 ;
        RECT 707.300 10.575 707.670 10.855 ;
        RECT 707.295 10.195 707.675 10.575 ;
        RECT 707.300 9.915 707.670 10.195 ;
        RECT 707.295 9.535 707.675 9.915 ;
        RECT 707.300 9.255 707.670 9.535 ;
        RECT 707.295 8.875 707.675 9.255 ;
        RECT 710.120 9.185 710.560 59.185 ;
        RECT 710.150 8.875 710.530 9.185 ;
        RECT 710.910 9.175 711.290 59.195 ;
        RECT 711.940 55.495 712.310 59.195 ;
        RECT 711.935 55.115 712.315 55.495 ;
        RECT 711.940 54.835 712.310 55.115 ;
        RECT 711.935 54.455 712.315 54.835 ;
        RECT 711.940 54.175 712.310 54.455 ;
        RECT 711.935 53.795 712.315 54.175 ;
        RECT 711.940 53.515 712.310 53.795 ;
        RECT 711.935 53.135 712.315 53.515 ;
        RECT 711.940 52.855 712.310 53.135 ;
        RECT 711.935 52.475 712.315 52.855 ;
        RECT 711.940 52.195 712.310 52.475 ;
        RECT 711.935 51.815 712.315 52.195 ;
        RECT 711.940 51.535 712.310 51.815 ;
        RECT 711.935 51.155 712.315 51.535 ;
        RECT 711.940 50.875 712.310 51.155 ;
        RECT 711.935 50.495 712.315 50.875 ;
        RECT 711.940 18.495 712.310 50.495 ;
        RECT 711.935 18.115 712.315 18.495 ;
        RECT 711.940 17.835 712.310 18.115 ;
        RECT 711.935 17.455 712.315 17.835 ;
        RECT 711.940 17.175 712.310 17.455 ;
        RECT 711.935 16.795 712.315 17.175 ;
        RECT 711.940 16.515 712.310 16.795 ;
        RECT 711.935 16.135 712.315 16.515 ;
        RECT 711.940 15.855 712.310 16.135 ;
        RECT 711.935 15.475 712.315 15.855 ;
        RECT 711.940 15.195 712.310 15.475 ;
        RECT 711.935 14.815 712.315 15.195 ;
        RECT 711.940 14.535 712.310 14.815 ;
        RECT 711.935 14.155 712.315 14.535 ;
        RECT 711.940 13.875 712.310 14.155 ;
        RECT 711.935 13.495 712.315 13.875 ;
        RECT 711.940 13.215 712.310 13.495 ;
        RECT 711.935 12.835 712.315 13.215 ;
        RECT 711.940 12.555 712.310 12.835 ;
        RECT 711.935 12.175 712.315 12.555 ;
        RECT 711.940 11.895 712.310 12.175 ;
        RECT 711.935 11.515 712.315 11.895 ;
        RECT 711.940 11.235 712.310 11.515 ;
        RECT 711.935 10.855 712.315 11.235 ;
        RECT 711.940 10.575 712.310 10.855 ;
        RECT 711.935 10.195 712.315 10.575 ;
        RECT 711.940 9.915 712.310 10.195 ;
        RECT 711.935 9.535 712.315 9.915 ;
        RECT 711.940 9.255 712.310 9.535 ;
        RECT 711.935 8.875 712.315 9.255 ;
        RECT 714.760 9.185 715.200 59.185 ;
        RECT 714.790 8.875 715.170 9.185 ;
        RECT 715.550 9.175 715.930 59.195 ;
        RECT 716.580 55.495 716.950 59.195 ;
        RECT 716.575 55.115 716.955 55.495 ;
        RECT 716.580 54.835 716.950 55.115 ;
        RECT 716.575 54.455 716.955 54.835 ;
        RECT 716.580 54.175 716.950 54.455 ;
        RECT 716.575 53.795 716.955 54.175 ;
        RECT 716.580 53.515 716.950 53.795 ;
        RECT 716.575 53.135 716.955 53.515 ;
        RECT 716.580 52.855 716.950 53.135 ;
        RECT 716.575 52.475 716.955 52.855 ;
        RECT 716.580 52.195 716.950 52.475 ;
        RECT 716.575 51.815 716.955 52.195 ;
        RECT 716.580 51.535 716.950 51.815 ;
        RECT 716.575 51.155 716.955 51.535 ;
        RECT 716.580 50.875 716.950 51.155 ;
        RECT 716.575 50.495 716.955 50.875 ;
        RECT 716.580 18.495 716.950 50.495 ;
        RECT 716.575 18.115 716.955 18.495 ;
        RECT 716.580 17.835 716.950 18.115 ;
        RECT 716.575 17.455 716.955 17.835 ;
        RECT 716.580 17.175 716.950 17.455 ;
        RECT 716.575 16.795 716.955 17.175 ;
        RECT 716.580 16.515 716.950 16.795 ;
        RECT 716.575 16.135 716.955 16.515 ;
        RECT 716.580 15.855 716.950 16.135 ;
        RECT 716.575 15.475 716.955 15.855 ;
        RECT 716.580 15.195 716.950 15.475 ;
        RECT 716.575 14.815 716.955 15.195 ;
        RECT 716.580 14.535 716.950 14.815 ;
        RECT 716.575 14.155 716.955 14.535 ;
        RECT 716.580 13.875 716.950 14.155 ;
        RECT 716.575 13.495 716.955 13.875 ;
        RECT 716.580 13.215 716.950 13.495 ;
        RECT 716.575 12.835 716.955 13.215 ;
        RECT 716.580 12.555 716.950 12.835 ;
        RECT 716.575 12.175 716.955 12.555 ;
        RECT 716.580 11.895 716.950 12.175 ;
        RECT 716.575 11.515 716.955 11.895 ;
        RECT 716.580 11.235 716.950 11.515 ;
        RECT 716.575 10.855 716.955 11.235 ;
        RECT 716.580 10.575 716.950 10.855 ;
        RECT 716.575 10.195 716.955 10.575 ;
        RECT 716.580 9.915 716.950 10.195 ;
        RECT 716.575 9.535 716.955 9.915 ;
        RECT 716.580 9.255 716.950 9.535 ;
        RECT 716.575 8.875 716.955 9.255 ;
        RECT 0.500 4.580 2.740 5.180 ;
        RECT 0.870 3.690 1.210 4.580 ;
        RECT 2.010 3.695 2.350 4.580 ;
        RECT 3.490 4.030 3.860 4.550 ;
        RECT 4.610 4.030 4.990 8.470 ;
        RECT 5.340 4.580 20.930 5.180 ;
        RECT 5.340 4.040 5.780 4.580 ;
        RECT 4.170 3.740 4.550 3.800 ;
        RECT 3.455 3.420 4.550 3.740 ;
        RECT 6.615 3.720 6.845 4.580 ;
        RECT 3.455 3.410 4.540 3.420 ;
        RECT 0.870 1.260 1.210 2.960 ;
        RECT 2.010 1.260 2.350 2.950 ;
        RECT 4.270 2.820 5.270 3.150 ;
        RECT 4.580 2.760 4.960 2.820 ;
        RECT 7.080 2.680 7.405 3.680 ;
        RECT 7.635 3.330 7.965 4.350 ;
        RECT 8.855 3.720 9.085 4.580 ;
        RECT 9.320 3.330 9.645 3.680 ;
        RECT 7.635 3.065 9.645 3.330 ;
        RECT 0.500 0.660 2.740 1.260 ;
        RECT 3.820 0.610 4.190 2.530 ;
        RECT 4.840 1.260 5.220 2.530 ;
        RECT 5.570 1.260 6.010 2.520 ;
        RECT 6.715 1.260 6.945 2.350 ;
        RECT 7.635 1.490 7.965 3.065 ;
        RECT 9.320 2.680 9.645 3.065 ;
        RECT 8.955 1.260 9.185 2.350 ;
        RECT 9.875 1.490 10.205 4.350 ;
        RECT 11.095 3.930 11.325 4.580 ;
        RECT 12.245 3.660 12.475 4.350 ;
        RECT 13.365 3.930 13.595 4.580 ;
        RECT 12.245 3.405 13.530 3.660 ;
        RECT 11.480 2.760 13.000 3.175 ;
        RECT 13.230 2.520 13.530 3.405 ;
        RECT 11.095 1.260 11.325 2.240 ;
        RECT 12.070 2.200 13.530 2.520 ;
        RECT 14.455 2.300 14.685 4.080 ;
        RECT 14.915 3.250 15.430 4.230 ;
        RECT 15.795 4.015 16.025 4.580 ;
        RECT 16.540 3.280 17.165 4.305 ;
        RECT 14.915 2.690 15.800 3.250 ;
        RECT 16.180 2.300 16.465 3.050 ;
        RECT 12.070 1.490 12.520 2.200 ;
        RECT 14.455 2.065 16.465 2.300 ;
        RECT 13.365 1.260 13.595 1.950 ;
        RECT 14.455 1.490 14.840 2.065 ;
        RECT 15.740 1.260 16.080 1.750 ;
        RECT 16.695 1.500 17.165 3.280 ;
        RECT 17.815 2.300 18.045 4.080 ;
        RECT 18.275 3.250 18.790 4.230 ;
        RECT 19.155 4.015 19.385 4.580 ;
        RECT 19.900 3.280 20.525 4.305 ;
        RECT 21.680 4.030 22.050 4.550 ;
        RECT 22.800 4.030 23.180 8.470 ;
        RECT 23.530 4.580 36.880 5.180 ;
        RECT 23.530 4.040 23.970 4.580 ;
        RECT 22.360 3.740 22.740 3.800 ;
        RECT 21.645 3.420 22.740 3.740 ;
        RECT 24.805 3.720 25.035 4.580 ;
        RECT 21.645 3.410 22.730 3.420 ;
        RECT 18.275 2.690 19.160 3.250 ;
        RECT 19.540 2.300 19.825 3.050 ;
        RECT 17.815 2.065 19.825 2.300 ;
        RECT 17.815 1.490 18.200 2.065 ;
        RECT 19.100 1.260 19.440 1.750 ;
        RECT 20.055 1.500 20.525 3.280 ;
        RECT 22.460 2.820 23.460 3.150 ;
        RECT 22.770 2.760 23.150 2.820 ;
        RECT 25.270 2.680 25.595 3.680 ;
        RECT 25.825 3.330 26.155 4.350 ;
        RECT 27.045 3.720 27.275 4.580 ;
        RECT 27.510 3.330 27.835 3.680 ;
        RECT 25.825 3.065 27.835 3.330 ;
        RECT 4.840 0.660 20.930 1.260 ;
        RECT 4.840 0.610 5.220 0.660 ;
        RECT 5.570 0.620 6.010 0.660 ;
        RECT 22.010 0.610 22.380 2.530 ;
        RECT 23.030 1.260 23.410 2.530 ;
        RECT 23.760 1.260 24.200 2.520 ;
        RECT 24.905 1.260 25.135 2.350 ;
        RECT 25.825 1.490 26.155 3.065 ;
        RECT 27.510 2.680 27.835 3.065 ;
        RECT 27.145 1.260 27.375 2.350 ;
        RECT 28.065 1.490 28.395 4.350 ;
        RECT 29.285 3.930 29.515 4.580 ;
        RECT 30.435 3.660 30.665 4.350 ;
        RECT 31.555 3.930 31.785 4.580 ;
        RECT 30.435 3.405 31.720 3.660 ;
        RECT 29.670 2.760 31.190 3.175 ;
        RECT 31.420 2.520 31.720 3.405 ;
        RECT 29.285 1.260 29.515 2.240 ;
        RECT 30.260 2.200 31.720 2.520 ;
        RECT 32.645 2.300 32.875 4.080 ;
        RECT 33.105 3.250 33.620 4.230 ;
        RECT 33.985 4.015 34.215 4.580 ;
        RECT 34.730 3.280 35.355 4.305 ;
        RECT 36.150 3.695 36.490 4.580 ;
        RECT 37.630 4.030 38.000 4.550 ;
        RECT 38.750 4.030 39.130 8.470 ;
        RECT 39.480 4.580 51.710 5.180 ;
        RECT 39.480 4.040 39.920 4.580 ;
        RECT 38.310 3.740 38.690 3.800 ;
        RECT 37.595 3.420 38.690 3.740 ;
        RECT 40.755 3.720 40.985 4.580 ;
        RECT 37.595 3.410 38.680 3.420 ;
        RECT 33.105 2.690 33.990 3.250 ;
        RECT 34.370 2.300 34.655 3.050 ;
        RECT 30.260 1.490 30.710 2.200 ;
        RECT 32.645 2.065 34.655 2.300 ;
        RECT 31.555 1.260 31.785 1.950 ;
        RECT 32.645 1.490 33.030 2.065 ;
        RECT 33.930 1.260 34.270 1.750 ;
        RECT 34.885 1.500 35.355 3.280 ;
        RECT 36.150 1.260 36.490 2.950 ;
        RECT 38.410 2.820 39.410 3.150 ;
        RECT 38.720 2.760 39.100 2.820 ;
        RECT 41.220 2.680 41.545 3.680 ;
        RECT 41.775 3.330 42.105 4.350 ;
        RECT 42.995 3.720 43.225 4.580 ;
        RECT 43.460 3.330 43.785 3.680 ;
        RECT 41.775 3.065 43.785 3.330 ;
        RECT 23.030 0.660 36.880 1.260 ;
        RECT 23.030 0.610 23.410 0.660 ;
        RECT 23.760 0.620 24.200 0.660 ;
        RECT 37.960 0.610 38.330 2.530 ;
        RECT 38.980 1.260 39.360 2.530 ;
        RECT 39.710 1.260 40.150 2.520 ;
        RECT 40.855 1.260 41.085 2.350 ;
        RECT 41.775 1.490 42.105 3.065 ;
        RECT 43.460 2.680 43.785 3.065 ;
        RECT 43.095 1.260 43.325 2.350 ;
        RECT 44.015 1.490 44.345 4.350 ;
        RECT 45.235 3.930 45.465 4.580 ;
        RECT 46.385 3.660 46.615 4.350 ;
        RECT 47.505 3.930 47.735 4.580 ;
        RECT 46.385 3.405 47.670 3.660 ;
        RECT 45.620 2.760 47.140 3.175 ;
        RECT 47.370 2.520 47.670 3.405 ;
        RECT 45.235 1.260 45.465 2.240 ;
        RECT 46.210 2.200 47.670 2.520 ;
        RECT 48.595 2.300 48.825 4.080 ;
        RECT 49.055 3.250 49.570 4.230 ;
        RECT 49.935 4.015 50.165 4.580 ;
        RECT 50.680 3.280 51.305 4.305 ;
        RECT 52.460 4.030 52.830 4.550 ;
        RECT 53.580 4.030 53.960 8.470 ;
        RECT 54.310 4.580 71.020 5.180 ;
        RECT 54.310 4.040 54.750 4.580 ;
        RECT 53.140 3.740 53.520 3.800 ;
        RECT 52.425 3.420 53.520 3.740 ;
        RECT 55.585 3.720 55.815 4.580 ;
        RECT 52.425 3.410 53.510 3.420 ;
        RECT 49.055 2.690 49.940 3.250 ;
        RECT 50.320 2.300 50.605 3.050 ;
        RECT 46.210 1.490 46.660 2.200 ;
        RECT 48.595 2.065 50.605 2.300 ;
        RECT 47.505 1.260 47.735 1.950 ;
        RECT 48.595 1.490 48.980 2.065 ;
        RECT 49.880 1.260 50.220 1.750 ;
        RECT 50.835 1.500 51.305 3.280 ;
        RECT 53.240 2.820 54.240 3.150 ;
        RECT 53.550 2.760 53.930 2.820 ;
        RECT 56.050 2.680 56.375 3.680 ;
        RECT 56.605 3.330 56.935 4.350 ;
        RECT 57.825 3.720 58.055 4.580 ;
        RECT 58.290 3.330 58.615 3.680 ;
        RECT 56.605 3.065 58.615 3.330 ;
        RECT 38.980 0.660 51.710 1.260 ;
        RECT 38.980 0.610 39.360 0.660 ;
        RECT 39.710 0.620 40.150 0.660 ;
        RECT 52.790 0.610 53.160 2.530 ;
        RECT 53.810 1.260 54.190 2.530 ;
        RECT 54.540 1.260 54.980 2.520 ;
        RECT 55.685 1.260 55.915 2.350 ;
        RECT 56.605 1.490 56.935 3.065 ;
        RECT 58.290 2.680 58.615 3.065 ;
        RECT 57.925 1.260 58.155 2.350 ;
        RECT 58.845 1.490 59.175 4.350 ;
        RECT 60.065 3.930 60.295 4.580 ;
        RECT 61.215 3.660 61.445 4.350 ;
        RECT 62.335 3.930 62.565 4.580 ;
        RECT 61.215 3.405 62.500 3.660 ;
        RECT 60.450 2.760 61.970 3.175 ;
        RECT 62.200 2.520 62.500 3.405 ;
        RECT 60.065 1.260 60.295 2.240 ;
        RECT 61.040 2.200 62.500 2.520 ;
        RECT 63.425 2.300 63.655 4.080 ;
        RECT 63.885 3.250 64.400 4.230 ;
        RECT 64.765 4.015 64.995 4.580 ;
        RECT 65.510 3.280 66.135 4.305 ;
        RECT 63.885 2.690 64.770 3.250 ;
        RECT 65.150 2.300 65.435 3.050 ;
        RECT 61.040 1.490 61.490 2.200 ;
        RECT 63.425 2.065 65.435 2.300 ;
        RECT 62.335 1.260 62.565 1.950 ;
        RECT 63.425 1.490 63.810 2.065 ;
        RECT 64.710 1.260 65.050 1.750 ;
        RECT 65.665 1.500 66.135 3.280 ;
        RECT 66.785 2.300 67.015 4.080 ;
        RECT 67.245 3.250 67.760 4.230 ;
        RECT 68.125 4.015 68.355 4.580 ;
        RECT 68.870 3.280 69.495 4.305 ;
        RECT 70.290 3.695 70.630 4.580 ;
        RECT 71.770 4.030 72.140 4.550 ;
        RECT 72.890 4.030 73.270 8.470 ;
        RECT 73.620 4.580 85.850 5.180 ;
        RECT 73.620 4.040 74.060 4.580 ;
        RECT 72.450 3.740 72.830 3.800 ;
        RECT 71.735 3.420 72.830 3.740 ;
        RECT 74.895 3.720 75.125 4.580 ;
        RECT 71.735 3.410 72.820 3.420 ;
        RECT 67.245 2.690 68.130 3.250 ;
        RECT 68.510 2.300 68.795 3.050 ;
        RECT 66.785 2.065 68.795 2.300 ;
        RECT 66.785 1.490 67.170 2.065 ;
        RECT 68.070 1.260 68.410 1.750 ;
        RECT 69.025 1.500 69.495 3.280 ;
        RECT 70.290 1.260 70.630 2.950 ;
        RECT 72.550 2.820 73.550 3.150 ;
        RECT 72.860 2.760 73.240 2.820 ;
        RECT 75.360 2.680 75.685 3.680 ;
        RECT 75.915 3.330 76.245 4.350 ;
        RECT 77.135 3.720 77.365 4.580 ;
        RECT 77.600 3.330 77.925 3.680 ;
        RECT 75.915 3.065 77.925 3.330 ;
        RECT 53.810 0.660 71.020 1.260 ;
        RECT 53.810 0.610 54.190 0.660 ;
        RECT 54.540 0.620 54.980 0.660 ;
        RECT 72.100 0.610 72.470 2.530 ;
        RECT 73.120 1.260 73.500 2.530 ;
        RECT 73.850 1.260 74.290 2.520 ;
        RECT 74.995 1.260 75.225 2.350 ;
        RECT 75.915 1.490 76.245 3.065 ;
        RECT 77.600 2.680 77.925 3.065 ;
        RECT 77.235 1.260 77.465 2.350 ;
        RECT 78.155 1.490 78.485 4.350 ;
        RECT 79.375 3.930 79.605 4.580 ;
        RECT 80.525 3.660 80.755 4.350 ;
        RECT 81.645 3.930 81.875 4.580 ;
        RECT 80.525 3.405 81.810 3.660 ;
        RECT 79.760 2.760 81.280 3.175 ;
        RECT 81.510 2.520 81.810 3.405 ;
        RECT 79.375 1.260 79.605 2.240 ;
        RECT 80.350 2.200 81.810 2.520 ;
        RECT 82.735 2.300 82.965 4.080 ;
        RECT 83.195 3.250 83.710 4.230 ;
        RECT 84.075 4.015 84.305 4.580 ;
        RECT 84.820 3.280 85.445 4.305 ;
        RECT 86.600 4.030 86.970 4.550 ;
        RECT 87.720 4.030 88.100 8.470 ;
        RECT 88.450 4.580 105.160 5.180 ;
        RECT 88.450 4.040 88.890 4.580 ;
        RECT 87.280 3.740 87.660 3.800 ;
        RECT 86.565 3.420 87.660 3.740 ;
        RECT 89.725 3.720 89.955 4.580 ;
        RECT 86.565 3.410 87.650 3.420 ;
        RECT 83.195 2.690 84.080 3.250 ;
        RECT 84.460 2.300 84.745 3.050 ;
        RECT 80.350 1.490 80.800 2.200 ;
        RECT 82.735 2.065 84.745 2.300 ;
        RECT 81.645 1.260 81.875 1.950 ;
        RECT 82.735 1.490 83.120 2.065 ;
        RECT 84.020 1.260 84.360 1.750 ;
        RECT 84.975 1.500 85.445 3.280 ;
        RECT 87.380 2.820 88.380 3.150 ;
        RECT 87.690 2.760 88.070 2.820 ;
        RECT 90.190 2.680 90.515 3.680 ;
        RECT 90.745 3.330 91.075 4.350 ;
        RECT 91.965 3.720 92.195 4.580 ;
        RECT 92.430 3.330 92.755 3.680 ;
        RECT 90.745 3.065 92.755 3.330 ;
        RECT 73.120 0.660 85.850 1.260 ;
        RECT 73.120 0.610 73.500 0.660 ;
        RECT 73.850 0.620 74.290 0.660 ;
        RECT 86.930 0.610 87.300 2.530 ;
        RECT 87.950 1.260 88.330 2.530 ;
        RECT 88.680 1.260 89.120 2.520 ;
        RECT 89.825 1.260 90.055 2.350 ;
        RECT 90.745 1.490 91.075 3.065 ;
        RECT 92.430 2.680 92.755 3.065 ;
        RECT 92.065 1.260 92.295 2.350 ;
        RECT 92.985 1.490 93.315 4.350 ;
        RECT 94.205 3.930 94.435 4.580 ;
        RECT 95.355 3.660 95.585 4.350 ;
        RECT 96.475 3.930 96.705 4.580 ;
        RECT 95.355 3.405 96.640 3.660 ;
        RECT 94.590 2.760 96.110 3.175 ;
        RECT 96.340 2.520 96.640 3.405 ;
        RECT 94.205 1.260 94.435 2.240 ;
        RECT 95.180 2.200 96.640 2.520 ;
        RECT 97.565 2.300 97.795 4.080 ;
        RECT 98.025 3.250 98.540 4.230 ;
        RECT 98.905 4.015 99.135 4.580 ;
        RECT 99.650 3.280 100.275 4.305 ;
        RECT 98.025 2.690 98.910 3.250 ;
        RECT 99.290 2.300 99.575 3.050 ;
        RECT 95.180 1.490 95.630 2.200 ;
        RECT 97.565 2.065 99.575 2.300 ;
        RECT 96.475 1.260 96.705 1.950 ;
        RECT 97.565 1.490 97.950 2.065 ;
        RECT 98.850 1.260 99.190 1.750 ;
        RECT 99.805 1.500 100.275 3.280 ;
        RECT 100.925 2.300 101.155 4.080 ;
        RECT 101.385 3.250 101.900 4.230 ;
        RECT 102.265 4.015 102.495 4.580 ;
        RECT 103.010 3.280 103.635 4.305 ;
        RECT 104.430 3.695 104.770 4.580 ;
        RECT 105.910 4.030 106.280 4.550 ;
        RECT 107.030 4.030 107.410 8.470 ;
        RECT 107.760 4.580 119.990 5.180 ;
        RECT 107.760 4.040 108.200 4.580 ;
        RECT 106.590 3.740 106.970 3.800 ;
        RECT 105.875 3.420 106.970 3.740 ;
        RECT 109.035 3.720 109.265 4.580 ;
        RECT 105.875 3.410 106.960 3.420 ;
        RECT 101.385 2.690 102.270 3.250 ;
        RECT 102.650 2.300 102.935 3.050 ;
        RECT 100.925 2.065 102.935 2.300 ;
        RECT 100.925 1.490 101.310 2.065 ;
        RECT 102.210 1.260 102.550 1.750 ;
        RECT 103.165 1.500 103.635 3.280 ;
        RECT 104.430 1.260 104.770 2.950 ;
        RECT 106.690 2.820 107.690 3.150 ;
        RECT 107.000 2.760 107.380 2.820 ;
        RECT 109.500 2.680 109.825 3.680 ;
        RECT 110.055 3.330 110.385 4.350 ;
        RECT 111.275 3.720 111.505 4.580 ;
        RECT 111.740 3.330 112.065 3.680 ;
        RECT 110.055 3.065 112.065 3.330 ;
        RECT 87.950 0.660 105.160 1.260 ;
        RECT 87.950 0.610 88.330 0.660 ;
        RECT 88.680 0.620 89.120 0.660 ;
        RECT 106.240 0.610 106.610 2.530 ;
        RECT 107.260 1.260 107.640 2.530 ;
        RECT 107.990 1.260 108.430 2.520 ;
        RECT 109.135 1.260 109.365 2.350 ;
        RECT 110.055 1.490 110.385 3.065 ;
        RECT 111.740 2.680 112.065 3.065 ;
        RECT 111.375 1.260 111.605 2.350 ;
        RECT 112.295 1.490 112.625 4.350 ;
        RECT 113.515 3.930 113.745 4.580 ;
        RECT 114.665 3.660 114.895 4.350 ;
        RECT 115.785 3.930 116.015 4.580 ;
        RECT 114.665 3.405 115.950 3.660 ;
        RECT 113.900 2.760 115.420 3.175 ;
        RECT 115.650 2.520 115.950 3.405 ;
        RECT 113.515 1.260 113.745 2.240 ;
        RECT 114.490 2.200 115.950 2.520 ;
        RECT 116.875 2.300 117.105 4.080 ;
        RECT 117.335 3.250 117.850 4.230 ;
        RECT 118.215 4.015 118.445 4.580 ;
        RECT 118.960 3.280 119.585 4.305 ;
        RECT 120.740 4.030 121.110 4.550 ;
        RECT 121.860 4.030 122.240 8.470 ;
        RECT 122.590 4.580 680.260 5.180 ;
        RECT 122.590 4.040 123.030 4.580 ;
        RECT 121.420 3.740 121.800 3.800 ;
        RECT 120.705 3.420 121.800 3.740 ;
        RECT 123.865 3.720 124.095 4.580 ;
        RECT 120.705 3.410 121.790 3.420 ;
        RECT 117.335 2.690 118.220 3.250 ;
        RECT 118.600 2.300 118.885 3.050 ;
        RECT 114.490 1.490 114.940 2.200 ;
        RECT 116.875 2.065 118.885 2.300 ;
        RECT 115.785 1.260 116.015 1.950 ;
        RECT 116.875 1.490 117.260 2.065 ;
        RECT 118.160 1.260 118.500 1.750 ;
        RECT 119.115 1.500 119.585 3.280 ;
        RECT 121.520 2.820 122.520 3.150 ;
        RECT 121.830 2.760 122.210 2.820 ;
        RECT 124.330 2.680 124.655 3.680 ;
        RECT 124.885 3.330 125.215 4.350 ;
        RECT 126.105 3.720 126.335 4.580 ;
        RECT 126.570 3.330 126.895 3.680 ;
        RECT 124.885 3.065 126.895 3.330 ;
        RECT 107.260 0.660 119.990 1.260 ;
        RECT 107.260 0.610 107.640 0.660 ;
        RECT 107.990 0.620 108.430 0.660 ;
        RECT 121.070 0.610 121.440 2.530 ;
        RECT 122.090 1.260 122.470 2.530 ;
        RECT 122.820 1.260 123.260 2.520 ;
        RECT 123.965 1.260 124.195 2.350 ;
        RECT 124.885 1.490 125.215 3.065 ;
        RECT 126.570 2.680 126.895 3.065 ;
        RECT 126.205 1.260 126.435 2.350 ;
        RECT 127.125 1.490 127.455 4.350 ;
        RECT 128.345 3.930 128.575 4.580 ;
        RECT 129.495 3.660 129.725 4.350 ;
        RECT 130.615 3.930 130.845 4.580 ;
        RECT 129.495 3.405 130.780 3.660 ;
        RECT 128.730 2.760 130.250 3.175 ;
        RECT 130.480 2.520 130.780 3.405 ;
        RECT 128.345 1.260 128.575 2.240 ;
        RECT 129.320 2.200 130.780 2.520 ;
        RECT 131.705 2.300 131.935 4.080 ;
        RECT 132.165 3.250 132.680 4.230 ;
        RECT 133.045 4.015 133.275 4.580 ;
        RECT 133.790 3.280 134.415 4.305 ;
        RECT 135.210 3.695 135.550 4.580 ;
        RECT 136.185 3.785 136.415 4.580 ;
        RECT 132.165 2.690 133.050 3.250 ;
        RECT 133.430 2.300 133.715 3.050 ;
        RECT 129.320 1.490 129.770 2.200 ;
        RECT 131.705 2.065 133.715 2.300 ;
        RECT 130.615 1.260 130.845 1.950 ;
        RECT 131.705 1.490 132.090 2.065 ;
        RECT 132.990 1.260 133.330 1.750 ;
        RECT 133.945 1.500 134.415 3.280 ;
        RECT 136.185 3.325 137.460 3.555 ;
        RECT 135.210 1.260 135.550 2.950 ;
        RECT 136.185 1.490 136.415 3.325 ;
        RECT 137.705 2.920 137.935 4.350 ;
        RECT 138.425 3.785 138.655 4.580 ;
        RECT 136.670 2.690 137.935 2.920 ;
        RECT 138.425 3.325 139.700 3.555 ;
        RECT 137.705 1.260 137.935 2.390 ;
        RECT 138.425 1.490 138.655 3.325 ;
        RECT 139.945 2.920 140.175 4.350 ;
        RECT 138.910 2.690 140.175 2.920 ;
        RECT 139.945 1.260 140.175 2.390 ;
        RECT 140.665 2.300 140.895 4.080 ;
        RECT 141.125 3.250 141.640 4.230 ;
        RECT 142.005 4.015 142.235 4.580 ;
        RECT 142.750 3.280 143.375 4.305 ;
        RECT 144.025 3.785 144.255 4.580 ;
        RECT 141.125 2.690 142.010 3.250 ;
        RECT 142.390 2.300 142.675 3.050 ;
        RECT 140.665 2.065 142.675 2.300 ;
        RECT 140.665 1.490 141.050 2.065 ;
        RECT 141.950 1.260 142.290 1.750 ;
        RECT 142.905 1.500 143.375 3.280 ;
        RECT 144.025 3.325 145.300 3.555 ;
        RECT 144.025 1.490 144.255 3.325 ;
        RECT 145.545 2.920 145.775 4.350 ;
        RECT 146.265 3.785 146.495 4.580 ;
        RECT 144.510 2.690 145.775 2.920 ;
        RECT 146.265 3.325 147.540 3.555 ;
        RECT 145.545 1.260 145.775 2.390 ;
        RECT 146.265 1.490 146.495 3.325 ;
        RECT 147.785 2.920 148.015 4.350 ;
        RECT 148.505 3.785 148.735 4.580 ;
        RECT 146.750 2.690 148.015 2.920 ;
        RECT 148.505 3.325 149.780 3.555 ;
        RECT 147.785 1.260 148.015 2.390 ;
        RECT 148.505 1.490 148.735 3.325 ;
        RECT 150.025 2.920 150.255 4.350 ;
        RECT 150.745 3.785 150.975 4.580 ;
        RECT 148.990 2.690 150.255 2.920 ;
        RECT 150.745 3.325 152.020 3.555 ;
        RECT 150.025 1.260 150.255 2.390 ;
        RECT 150.745 1.490 150.975 3.325 ;
        RECT 152.265 2.920 152.495 4.350 ;
        RECT 152.985 3.785 153.215 4.580 ;
        RECT 151.230 2.690 152.495 2.920 ;
        RECT 152.985 3.325 154.260 3.555 ;
        RECT 152.265 1.260 152.495 2.390 ;
        RECT 152.985 1.490 153.215 3.325 ;
        RECT 154.505 2.920 154.735 4.350 ;
        RECT 155.370 3.695 155.710 4.580 ;
        RECT 156.345 3.785 156.575 4.580 ;
        RECT 156.345 3.325 157.620 3.555 ;
        RECT 153.470 2.690 154.735 2.920 ;
        RECT 154.505 1.260 154.735 2.390 ;
        RECT 155.370 1.260 155.710 2.950 ;
        RECT 156.345 1.490 156.575 3.325 ;
        RECT 157.865 2.920 158.095 4.350 ;
        RECT 158.585 3.785 158.815 4.580 ;
        RECT 156.830 2.690 158.095 2.920 ;
        RECT 158.585 3.325 159.860 3.555 ;
        RECT 157.865 1.260 158.095 2.390 ;
        RECT 158.585 1.490 158.815 3.325 ;
        RECT 160.105 2.920 160.335 4.350 ;
        RECT 160.825 3.785 161.055 4.580 ;
        RECT 159.070 2.690 160.335 2.920 ;
        RECT 160.825 3.325 162.100 3.555 ;
        RECT 160.105 1.260 160.335 2.390 ;
        RECT 160.825 1.490 161.055 3.325 ;
        RECT 162.345 2.920 162.575 4.350 ;
        RECT 163.065 3.785 163.295 4.580 ;
        RECT 161.310 2.690 162.575 2.920 ;
        RECT 163.065 3.325 164.340 3.555 ;
        RECT 162.345 1.260 162.575 2.390 ;
        RECT 163.065 1.490 163.295 3.325 ;
        RECT 164.585 2.920 164.815 4.350 ;
        RECT 165.305 3.785 165.535 4.580 ;
        RECT 163.550 2.690 164.815 2.920 ;
        RECT 165.305 3.325 166.580 3.555 ;
        RECT 164.585 1.260 164.815 2.390 ;
        RECT 165.305 1.490 165.535 3.325 ;
        RECT 166.825 2.920 167.055 4.350 ;
        RECT 167.545 3.785 167.775 4.580 ;
        RECT 165.790 2.690 167.055 2.920 ;
        RECT 167.545 3.325 168.820 3.555 ;
        RECT 166.825 1.260 167.055 2.390 ;
        RECT 167.545 1.490 167.775 3.325 ;
        RECT 169.065 2.920 169.295 4.350 ;
        RECT 169.785 3.785 170.015 4.580 ;
        RECT 168.030 2.690 169.295 2.920 ;
        RECT 169.785 3.325 171.060 3.555 ;
        RECT 169.065 1.260 169.295 2.390 ;
        RECT 169.785 1.490 170.015 3.325 ;
        RECT 171.305 2.920 171.535 4.350 ;
        RECT 172.025 3.785 172.255 4.580 ;
        RECT 170.270 2.690 171.535 2.920 ;
        RECT 172.025 3.325 173.300 3.555 ;
        RECT 171.305 1.260 171.535 2.390 ;
        RECT 172.025 1.490 172.255 3.325 ;
        RECT 173.545 2.920 173.775 4.350 ;
        RECT 174.265 3.785 174.495 4.580 ;
        RECT 172.510 2.690 173.775 2.920 ;
        RECT 174.265 3.325 175.540 3.555 ;
        RECT 173.545 1.260 173.775 2.390 ;
        RECT 174.265 1.490 174.495 3.325 ;
        RECT 175.785 2.920 176.015 4.350 ;
        RECT 176.650 3.695 176.990 4.580 ;
        RECT 177.625 3.785 177.855 4.580 ;
        RECT 177.625 3.325 178.900 3.555 ;
        RECT 174.750 2.690 176.015 2.920 ;
        RECT 175.785 1.260 176.015 2.390 ;
        RECT 176.650 1.260 176.990 2.950 ;
        RECT 177.625 1.490 177.855 3.325 ;
        RECT 179.145 2.920 179.375 4.350 ;
        RECT 179.865 3.785 180.095 4.580 ;
        RECT 178.110 2.690 179.375 2.920 ;
        RECT 179.865 3.325 181.140 3.555 ;
        RECT 179.145 1.260 179.375 2.390 ;
        RECT 179.865 1.490 180.095 3.325 ;
        RECT 181.385 2.920 181.615 4.350 ;
        RECT 180.350 2.690 181.615 2.920 ;
        RECT 181.385 1.260 181.615 2.390 ;
        RECT 182.105 2.300 182.335 4.080 ;
        RECT 182.565 3.250 183.080 4.230 ;
        RECT 183.445 4.015 183.675 4.580 ;
        RECT 184.190 3.280 184.815 4.305 ;
        RECT 185.465 3.785 185.695 4.580 ;
        RECT 182.565 2.690 183.450 3.250 ;
        RECT 183.830 2.300 184.115 3.050 ;
        RECT 182.105 2.065 184.115 2.300 ;
        RECT 182.105 1.490 182.490 2.065 ;
        RECT 183.390 1.260 183.730 1.750 ;
        RECT 184.345 1.500 184.815 3.280 ;
        RECT 185.465 3.325 186.740 3.555 ;
        RECT 185.465 1.490 185.695 3.325 ;
        RECT 186.985 2.920 187.215 4.350 ;
        RECT 187.705 3.785 187.935 4.580 ;
        RECT 185.950 2.690 187.215 2.920 ;
        RECT 187.705 3.325 188.980 3.555 ;
        RECT 186.985 1.260 187.215 2.390 ;
        RECT 187.705 1.490 187.935 3.325 ;
        RECT 189.225 2.920 189.455 4.350 ;
        RECT 189.945 3.785 190.175 4.580 ;
        RECT 188.190 2.690 189.455 2.920 ;
        RECT 189.945 3.325 191.220 3.555 ;
        RECT 189.225 1.260 189.455 2.390 ;
        RECT 189.945 1.490 190.175 3.325 ;
        RECT 191.465 2.920 191.695 4.350 ;
        RECT 192.185 3.785 192.415 4.580 ;
        RECT 190.430 2.690 191.695 2.920 ;
        RECT 192.185 3.325 193.460 3.555 ;
        RECT 191.465 1.260 191.695 2.390 ;
        RECT 192.185 1.490 192.415 3.325 ;
        RECT 193.705 2.920 193.935 4.350 ;
        RECT 194.425 3.785 194.655 4.580 ;
        RECT 192.670 2.690 193.935 2.920 ;
        RECT 194.425 3.325 195.700 3.555 ;
        RECT 193.705 1.260 193.935 2.390 ;
        RECT 194.425 1.490 194.655 3.325 ;
        RECT 195.945 2.920 196.175 4.350 ;
        RECT 196.810 3.695 197.150 4.580 ;
        RECT 197.785 3.785 198.015 4.580 ;
        RECT 197.785 3.325 199.060 3.555 ;
        RECT 194.910 2.690 196.175 2.920 ;
        RECT 195.945 1.260 196.175 2.390 ;
        RECT 196.810 1.260 197.150 2.950 ;
        RECT 197.785 1.490 198.015 3.325 ;
        RECT 199.305 2.920 199.535 4.350 ;
        RECT 200.025 3.785 200.255 4.580 ;
        RECT 198.270 2.690 199.535 2.920 ;
        RECT 200.025 3.325 201.300 3.555 ;
        RECT 199.305 1.260 199.535 2.390 ;
        RECT 200.025 1.490 200.255 3.325 ;
        RECT 201.545 2.920 201.775 4.350 ;
        RECT 202.265 3.785 202.495 4.580 ;
        RECT 200.510 2.690 201.775 2.920 ;
        RECT 202.265 3.325 203.540 3.555 ;
        RECT 201.545 1.260 201.775 2.390 ;
        RECT 202.265 1.490 202.495 3.325 ;
        RECT 203.785 2.920 204.015 4.350 ;
        RECT 204.505 3.785 204.735 4.580 ;
        RECT 202.750 2.690 204.015 2.920 ;
        RECT 204.505 3.325 205.780 3.555 ;
        RECT 203.785 1.260 204.015 2.390 ;
        RECT 204.505 1.490 204.735 3.325 ;
        RECT 206.025 2.920 206.255 4.350 ;
        RECT 206.745 3.785 206.975 4.580 ;
        RECT 204.990 2.690 206.255 2.920 ;
        RECT 206.745 3.325 208.020 3.555 ;
        RECT 206.025 1.260 206.255 2.390 ;
        RECT 206.745 1.490 206.975 3.325 ;
        RECT 208.265 2.920 208.495 4.350 ;
        RECT 208.985 3.785 209.215 4.580 ;
        RECT 207.230 2.690 208.495 2.920 ;
        RECT 208.985 3.325 210.260 3.555 ;
        RECT 208.265 1.260 208.495 2.390 ;
        RECT 208.985 1.490 209.215 3.325 ;
        RECT 210.505 2.920 210.735 4.350 ;
        RECT 211.225 3.785 211.455 4.580 ;
        RECT 209.470 2.690 210.735 2.920 ;
        RECT 211.225 3.325 212.500 3.555 ;
        RECT 210.505 1.260 210.735 2.390 ;
        RECT 211.225 1.490 211.455 3.325 ;
        RECT 212.745 2.920 212.975 4.350 ;
        RECT 213.465 3.785 213.695 4.580 ;
        RECT 211.710 2.690 212.975 2.920 ;
        RECT 213.465 3.325 214.740 3.555 ;
        RECT 212.745 1.260 212.975 2.390 ;
        RECT 213.465 1.490 213.695 3.325 ;
        RECT 214.985 2.920 215.215 4.350 ;
        RECT 215.705 3.785 215.935 4.580 ;
        RECT 213.950 2.690 215.215 2.920 ;
        RECT 215.705 3.325 216.980 3.555 ;
        RECT 214.985 1.260 215.215 2.390 ;
        RECT 215.705 1.490 215.935 3.325 ;
        RECT 217.225 2.920 217.455 4.350 ;
        RECT 218.090 3.695 218.430 4.580 ;
        RECT 219.065 3.785 219.295 4.580 ;
        RECT 219.065 3.325 220.340 3.555 ;
        RECT 216.190 2.690 217.455 2.920 ;
        RECT 217.225 1.260 217.455 2.390 ;
        RECT 218.090 1.260 218.430 2.950 ;
        RECT 219.065 1.490 219.295 3.325 ;
        RECT 220.585 2.920 220.815 4.350 ;
        RECT 221.305 3.785 221.535 4.580 ;
        RECT 219.550 2.690 220.815 2.920 ;
        RECT 221.305 3.325 222.580 3.555 ;
        RECT 220.585 1.260 220.815 2.390 ;
        RECT 221.305 1.490 221.535 3.325 ;
        RECT 222.825 2.920 223.055 4.350 ;
        RECT 223.545 3.785 223.775 4.580 ;
        RECT 221.790 2.690 223.055 2.920 ;
        RECT 223.545 3.325 224.820 3.555 ;
        RECT 222.825 1.260 223.055 2.390 ;
        RECT 223.545 1.490 223.775 3.325 ;
        RECT 225.065 2.920 225.295 4.350 ;
        RECT 224.030 2.690 225.295 2.920 ;
        RECT 225.065 1.260 225.295 2.390 ;
        RECT 225.785 2.300 226.015 4.080 ;
        RECT 226.245 3.250 226.760 4.230 ;
        RECT 227.125 4.015 227.355 4.580 ;
        RECT 227.870 3.280 228.495 4.305 ;
        RECT 229.145 3.785 229.375 4.580 ;
        RECT 226.245 2.690 227.130 3.250 ;
        RECT 227.510 2.300 227.795 3.050 ;
        RECT 225.785 2.065 227.795 2.300 ;
        RECT 225.785 1.490 226.170 2.065 ;
        RECT 227.070 1.260 227.410 1.750 ;
        RECT 228.025 1.500 228.495 3.280 ;
        RECT 229.145 3.325 230.420 3.555 ;
        RECT 229.145 1.490 229.375 3.325 ;
        RECT 230.665 2.920 230.895 4.350 ;
        RECT 231.385 3.785 231.615 4.580 ;
        RECT 229.630 2.690 230.895 2.920 ;
        RECT 231.385 3.325 232.660 3.555 ;
        RECT 230.665 1.260 230.895 2.390 ;
        RECT 231.385 1.490 231.615 3.325 ;
        RECT 232.905 2.920 233.135 4.350 ;
        RECT 233.625 3.785 233.855 4.580 ;
        RECT 231.870 2.690 233.135 2.920 ;
        RECT 233.625 3.325 234.900 3.555 ;
        RECT 232.905 1.260 233.135 2.390 ;
        RECT 233.625 1.490 233.855 3.325 ;
        RECT 235.145 2.920 235.375 4.350 ;
        RECT 235.865 3.785 236.095 4.580 ;
        RECT 234.110 2.690 235.375 2.920 ;
        RECT 235.865 3.325 237.140 3.555 ;
        RECT 235.145 1.260 235.375 2.390 ;
        RECT 235.865 1.490 236.095 3.325 ;
        RECT 237.385 2.920 237.615 4.350 ;
        RECT 238.250 3.695 238.590 4.580 ;
        RECT 239.225 3.785 239.455 4.580 ;
        RECT 239.225 3.325 240.500 3.555 ;
        RECT 236.350 2.690 237.615 2.920 ;
        RECT 237.385 1.260 237.615 2.390 ;
        RECT 238.250 1.260 238.590 2.950 ;
        RECT 239.225 1.490 239.455 3.325 ;
        RECT 240.745 2.920 240.975 4.350 ;
        RECT 241.465 3.785 241.695 4.580 ;
        RECT 239.710 2.690 240.975 2.920 ;
        RECT 241.465 3.325 242.740 3.555 ;
        RECT 240.745 1.260 240.975 2.390 ;
        RECT 241.465 1.490 241.695 3.325 ;
        RECT 242.985 2.920 243.215 4.350 ;
        RECT 243.705 3.785 243.935 4.580 ;
        RECT 241.950 2.690 243.215 2.920 ;
        RECT 243.705 3.325 244.980 3.555 ;
        RECT 242.985 1.260 243.215 2.390 ;
        RECT 243.705 1.490 243.935 3.325 ;
        RECT 245.225 2.920 245.455 4.350 ;
        RECT 245.945 3.785 246.175 4.580 ;
        RECT 244.190 2.690 245.455 2.920 ;
        RECT 245.945 3.325 247.220 3.555 ;
        RECT 245.225 1.260 245.455 2.390 ;
        RECT 245.945 1.490 246.175 3.325 ;
        RECT 247.465 2.920 247.695 4.350 ;
        RECT 248.185 3.785 248.415 4.580 ;
        RECT 246.430 2.690 247.695 2.920 ;
        RECT 248.185 3.325 249.460 3.555 ;
        RECT 247.465 1.260 247.695 2.390 ;
        RECT 248.185 1.490 248.415 3.325 ;
        RECT 249.705 2.920 249.935 4.350 ;
        RECT 250.425 3.785 250.655 4.580 ;
        RECT 248.670 2.690 249.935 2.920 ;
        RECT 250.425 3.325 251.700 3.555 ;
        RECT 249.705 1.260 249.935 2.390 ;
        RECT 250.425 1.490 250.655 3.325 ;
        RECT 251.945 2.920 252.175 4.350 ;
        RECT 252.665 3.785 252.895 4.580 ;
        RECT 250.910 2.690 252.175 2.920 ;
        RECT 252.665 3.325 253.940 3.555 ;
        RECT 251.945 1.260 252.175 2.390 ;
        RECT 252.665 1.490 252.895 3.325 ;
        RECT 254.185 2.920 254.415 4.350 ;
        RECT 254.905 3.785 255.135 4.580 ;
        RECT 253.150 2.690 254.415 2.920 ;
        RECT 254.905 3.325 256.180 3.555 ;
        RECT 254.185 1.260 254.415 2.390 ;
        RECT 254.905 1.490 255.135 3.325 ;
        RECT 256.425 2.920 256.655 4.350 ;
        RECT 257.145 3.785 257.375 4.580 ;
        RECT 255.390 2.690 256.655 2.920 ;
        RECT 257.145 3.325 258.420 3.555 ;
        RECT 256.425 1.260 256.655 2.390 ;
        RECT 257.145 1.490 257.375 3.325 ;
        RECT 258.665 2.920 258.895 4.350 ;
        RECT 259.530 3.695 259.870 4.580 ;
        RECT 260.505 3.785 260.735 4.580 ;
        RECT 260.505 3.325 261.780 3.555 ;
        RECT 257.630 2.690 258.895 2.920 ;
        RECT 258.665 1.260 258.895 2.390 ;
        RECT 259.530 1.260 259.870 2.950 ;
        RECT 260.505 1.490 260.735 3.325 ;
        RECT 262.025 2.920 262.255 4.350 ;
        RECT 262.745 3.785 262.975 4.580 ;
        RECT 260.990 2.690 262.255 2.920 ;
        RECT 262.745 3.325 264.020 3.555 ;
        RECT 262.025 1.260 262.255 2.390 ;
        RECT 262.745 1.490 262.975 3.325 ;
        RECT 264.265 2.920 264.495 4.350 ;
        RECT 264.985 3.785 265.215 4.580 ;
        RECT 263.230 2.690 264.495 2.920 ;
        RECT 264.985 3.325 266.260 3.555 ;
        RECT 264.265 1.260 264.495 2.390 ;
        RECT 264.985 1.490 265.215 3.325 ;
        RECT 266.505 2.920 266.735 4.350 ;
        RECT 265.470 2.690 266.735 2.920 ;
        RECT 266.505 1.260 266.735 2.390 ;
        RECT 267.225 2.300 267.455 4.080 ;
        RECT 267.685 3.250 268.200 4.230 ;
        RECT 268.565 4.015 268.795 4.580 ;
        RECT 269.310 3.280 269.935 4.305 ;
        RECT 270.585 3.785 270.815 4.580 ;
        RECT 267.685 2.690 268.570 3.250 ;
        RECT 268.950 2.300 269.235 3.050 ;
        RECT 267.225 2.065 269.235 2.300 ;
        RECT 267.225 1.490 267.610 2.065 ;
        RECT 268.510 1.260 268.850 1.750 ;
        RECT 269.465 1.500 269.935 3.280 ;
        RECT 270.585 3.325 271.860 3.555 ;
        RECT 270.585 1.490 270.815 3.325 ;
        RECT 272.105 2.920 272.335 4.350 ;
        RECT 272.825 3.785 273.055 4.580 ;
        RECT 271.070 2.690 272.335 2.920 ;
        RECT 272.825 3.325 274.100 3.555 ;
        RECT 272.105 1.260 272.335 2.390 ;
        RECT 272.825 1.490 273.055 3.325 ;
        RECT 274.345 2.920 274.575 4.350 ;
        RECT 275.065 3.785 275.295 4.580 ;
        RECT 273.310 2.690 274.575 2.920 ;
        RECT 275.065 3.325 276.340 3.555 ;
        RECT 274.345 1.260 274.575 2.390 ;
        RECT 275.065 1.490 275.295 3.325 ;
        RECT 276.585 2.920 276.815 4.350 ;
        RECT 277.305 3.785 277.535 4.580 ;
        RECT 275.550 2.690 276.815 2.920 ;
        RECT 277.305 3.325 278.580 3.555 ;
        RECT 276.585 1.260 276.815 2.390 ;
        RECT 277.305 1.490 277.535 3.325 ;
        RECT 278.825 2.920 279.055 4.350 ;
        RECT 279.690 3.695 280.030 4.580 ;
        RECT 280.665 3.785 280.895 4.580 ;
        RECT 280.665 3.325 281.940 3.555 ;
        RECT 277.790 2.690 279.055 2.920 ;
        RECT 278.825 1.260 279.055 2.390 ;
        RECT 279.690 1.260 280.030 2.950 ;
        RECT 280.665 1.490 280.895 3.325 ;
        RECT 282.185 2.920 282.415 4.350 ;
        RECT 282.905 3.785 283.135 4.580 ;
        RECT 281.150 2.690 282.415 2.920 ;
        RECT 282.905 3.325 284.180 3.555 ;
        RECT 282.185 1.260 282.415 2.390 ;
        RECT 282.905 1.490 283.135 3.325 ;
        RECT 284.425 2.920 284.655 4.350 ;
        RECT 285.145 3.785 285.375 4.580 ;
        RECT 283.390 2.690 284.655 2.920 ;
        RECT 285.145 3.325 286.420 3.555 ;
        RECT 284.425 1.260 284.655 2.390 ;
        RECT 285.145 1.490 285.375 3.325 ;
        RECT 286.665 2.920 286.895 4.350 ;
        RECT 287.385 3.785 287.615 4.580 ;
        RECT 285.630 2.690 286.895 2.920 ;
        RECT 287.385 3.325 288.660 3.555 ;
        RECT 286.665 1.260 286.895 2.390 ;
        RECT 287.385 1.490 287.615 3.325 ;
        RECT 288.905 2.920 289.135 4.350 ;
        RECT 289.625 3.785 289.855 4.580 ;
        RECT 287.870 2.690 289.135 2.920 ;
        RECT 289.625 3.325 290.900 3.555 ;
        RECT 288.905 1.260 289.135 2.390 ;
        RECT 289.625 1.490 289.855 3.325 ;
        RECT 291.145 2.920 291.375 4.350 ;
        RECT 291.865 3.785 292.095 4.580 ;
        RECT 290.110 2.690 291.375 2.920 ;
        RECT 291.865 3.325 293.140 3.555 ;
        RECT 291.145 1.260 291.375 2.390 ;
        RECT 291.865 1.490 292.095 3.325 ;
        RECT 293.385 2.920 293.615 4.350 ;
        RECT 294.105 3.785 294.335 4.580 ;
        RECT 292.350 2.690 293.615 2.920 ;
        RECT 294.105 3.325 295.380 3.555 ;
        RECT 293.385 1.260 293.615 2.390 ;
        RECT 294.105 1.490 294.335 3.325 ;
        RECT 295.625 2.920 295.855 4.350 ;
        RECT 296.345 3.785 296.575 4.580 ;
        RECT 294.590 2.690 295.855 2.920 ;
        RECT 296.345 3.325 297.620 3.555 ;
        RECT 295.625 1.260 295.855 2.390 ;
        RECT 296.345 1.490 296.575 3.325 ;
        RECT 297.865 2.920 298.095 4.350 ;
        RECT 298.585 3.785 298.815 4.580 ;
        RECT 296.830 2.690 298.095 2.920 ;
        RECT 298.585 3.325 299.860 3.555 ;
        RECT 297.865 1.260 298.095 2.390 ;
        RECT 298.585 1.490 298.815 3.325 ;
        RECT 300.105 2.920 300.335 4.350 ;
        RECT 300.970 3.695 301.310 4.580 ;
        RECT 301.945 3.785 302.175 4.580 ;
        RECT 301.945 3.325 303.220 3.555 ;
        RECT 299.070 2.690 300.335 2.920 ;
        RECT 300.105 1.260 300.335 2.390 ;
        RECT 300.970 1.260 301.310 2.950 ;
        RECT 301.945 1.490 302.175 3.325 ;
        RECT 303.465 2.920 303.695 4.350 ;
        RECT 304.185 3.785 304.415 4.580 ;
        RECT 302.430 2.690 303.695 2.920 ;
        RECT 304.185 3.325 305.460 3.555 ;
        RECT 303.465 1.260 303.695 2.390 ;
        RECT 304.185 1.490 304.415 3.325 ;
        RECT 305.705 2.920 305.935 4.350 ;
        RECT 306.425 3.785 306.655 4.580 ;
        RECT 304.670 2.690 305.935 2.920 ;
        RECT 306.425 3.325 307.700 3.555 ;
        RECT 305.705 1.260 305.935 2.390 ;
        RECT 306.425 1.490 306.655 3.325 ;
        RECT 307.945 2.920 308.175 4.350 ;
        RECT 308.665 3.785 308.895 4.580 ;
        RECT 306.910 2.690 308.175 2.920 ;
        RECT 308.665 3.325 309.940 3.555 ;
        RECT 307.945 1.260 308.175 2.390 ;
        RECT 308.665 1.490 308.895 3.325 ;
        RECT 310.185 2.920 310.415 4.350 ;
        RECT 309.150 2.690 310.415 2.920 ;
        RECT 310.185 1.260 310.415 2.390 ;
        RECT 310.905 2.300 311.135 4.080 ;
        RECT 311.365 3.250 311.880 4.230 ;
        RECT 312.245 4.015 312.475 4.580 ;
        RECT 312.990 3.280 313.615 4.305 ;
        RECT 314.265 3.785 314.495 4.580 ;
        RECT 311.365 2.690 312.250 3.250 ;
        RECT 312.630 2.300 312.915 3.050 ;
        RECT 310.905 2.065 312.915 2.300 ;
        RECT 310.905 1.490 311.290 2.065 ;
        RECT 312.190 1.260 312.530 1.750 ;
        RECT 313.145 1.500 313.615 3.280 ;
        RECT 314.265 3.325 315.540 3.555 ;
        RECT 314.265 1.490 314.495 3.325 ;
        RECT 315.785 2.920 316.015 4.350 ;
        RECT 316.505 3.785 316.735 4.580 ;
        RECT 314.750 2.690 316.015 2.920 ;
        RECT 316.505 3.325 317.780 3.555 ;
        RECT 315.785 1.260 316.015 2.390 ;
        RECT 316.505 1.490 316.735 3.325 ;
        RECT 318.025 2.920 318.255 4.350 ;
        RECT 318.745 3.785 318.975 4.580 ;
        RECT 316.990 2.690 318.255 2.920 ;
        RECT 318.745 3.325 320.020 3.555 ;
        RECT 318.025 1.260 318.255 2.390 ;
        RECT 318.745 1.490 318.975 3.325 ;
        RECT 320.265 2.920 320.495 4.350 ;
        RECT 321.130 3.695 321.470 4.580 ;
        RECT 322.105 3.785 322.335 4.580 ;
        RECT 322.105 3.325 323.380 3.555 ;
        RECT 319.230 2.690 320.495 2.920 ;
        RECT 320.265 1.260 320.495 2.390 ;
        RECT 321.130 1.260 321.470 2.950 ;
        RECT 322.105 1.490 322.335 3.325 ;
        RECT 323.625 2.920 323.855 4.350 ;
        RECT 324.345 3.785 324.575 4.580 ;
        RECT 322.590 2.690 323.855 2.920 ;
        RECT 324.345 3.325 325.620 3.555 ;
        RECT 323.625 1.260 323.855 2.390 ;
        RECT 324.345 1.490 324.575 3.325 ;
        RECT 325.865 2.920 326.095 4.350 ;
        RECT 326.585 3.785 326.815 4.580 ;
        RECT 324.830 2.690 326.095 2.920 ;
        RECT 326.585 3.325 327.860 3.555 ;
        RECT 325.865 1.260 326.095 2.390 ;
        RECT 326.585 1.490 326.815 3.325 ;
        RECT 328.105 2.920 328.335 4.350 ;
        RECT 328.825 3.785 329.055 4.580 ;
        RECT 327.070 2.690 328.335 2.920 ;
        RECT 328.825 3.325 330.100 3.555 ;
        RECT 328.105 1.260 328.335 2.390 ;
        RECT 328.825 1.490 329.055 3.325 ;
        RECT 330.345 2.920 330.575 4.350 ;
        RECT 331.065 3.785 331.295 4.580 ;
        RECT 329.310 2.690 330.575 2.920 ;
        RECT 331.065 3.325 332.340 3.555 ;
        RECT 330.345 1.260 330.575 2.390 ;
        RECT 331.065 1.490 331.295 3.325 ;
        RECT 332.585 2.920 332.815 4.350 ;
        RECT 333.305 3.785 333.535 4.580 ;
        RECT 331.550 2.690 332.815 2.920 ;
        RECT 333.305 3.325 334.580 3.555 ;
        RECT 332.585 1.260 332.815 2.390 ;
        RECT 333.305 1.490 333.535 3.325 ;
        RECT 334.825 2.920 335.055 4.350 ;
        RECT 335.545 3.785 335.775 4.580 ;
        RECT 333.790 2.690 335.055 2.920 ;
        RECT 335.545 3.325 336.820 3.555 ;
        RECT 334.825 1.260 335.055 2.390 ;
        RECT 335.545 1.490 335.775 3.325 ;
        RECT 337.065 2.920 337.295 4.350 ;
        RECT 337.785 3.785 338.015 4.580 ;
        RECT 336.030 2.690 337.295 2.920 ;
        RECT 337.785 3.325 339.060 3.555 ;
        RECT 337.065 1.260 337.295 2.390 ;
        RECT 337.785 1.490 338.015 3.325 ;
        RECT 339.305 2.920 339.535 4.350 ;
        RECT 340.025 3.785 340.255 4.580 ;
        RECT 338.270 2.690 339.535 2.920 ;
        RECT 340.025 3.325 341.300 3.555 ;
        RECT 339.305 1.260 339.535 2.390 ;
        RECT 340.025 1.490 340.255 3.325 ;
        RECT 341.545 2.920 341.775 4.350 ;
        RECT 342.410 3.695 342.750 4.580 ;
        RECT 343.385 3.785 343.615 4.580 ;
        RECT 343.385 3.325 344.660 3.555 ;
        RECT 340.510 2.690 341.775 2.920 ;
        RECT 341.545 1.260 341.775 2.390 ;
        RECT 342.410 1.260 342.750 2.950 ;
        RECT 343.385 1.490 343.615 3.325 ;
        RECT 344.905 2.920 345.135 4.350 ;
        RECT 345.625 3.785 345.855 4.580 ;
        RECT 343.870 2.690 345.135 2.920 ;
        RECT 345.625 3.325 346.900 3.555 ;
        RECT 344.905 1.260 345.135 2.390 ;
        RECT 345.625 1.490 345.855 3.325 ;
        RECT 347.145 2.920 347.375 4.350 ;
        RECT 347.865 3.785 348.095 4.580 ;
        RECT 346.110 2.690 347.375 2.920 ;
        RECT 347.865 3.325 349.140 3.555 ;
        RECT 347.145 1.260 347.375 2.390 ;
        RECT 347.865 1.490 348.095 3.325 ;
        RECT 349.385 2.920 349.615 4.350 ;
        RECT 350.105 3.785 350.335 4.580 ;
        RECT 348.350 2.690 349.615 2.920 ;
        RECT 350.105 3.325 351.380 3.555 ;
        RECT 349.385 1.260 349.615 2.390 ;
        RECT 350.105 1.490 350.335 3.325 ;
        RECT 351.625 2.920 351.855 4.350 ;
        RECT 350.590 2.690 351.855 2.920 ;
        RECT 351.625 1.260 351.855 2.390 ;
        RECT 352.345 2.300 352.575 4.080 ;
        RECT 352.805 3.250 353.320 4.230 ;
        RECT 353.685 4.015 353.915 4.580 ;
        RECT 354.430 3.280 355.055 4.305 ;
        RECT 355.705 3.785 355.935 4.580 ;
        RECT 352.805 2.690 353.690 3.250 ;
        RECT 354.070 2.300 354.355 3.050 ;
        RECT 352.345 2.065 354.355 2.300 ;
        RECT 352.345 1.490 352.730 2.065 ;
        RECT 353.630 1.260 353.970 1.750 ;
        RECT 354.585 1.500 355.055 3.280 ;
        RECT 355.705 3.325 356.980 3.555 ;
        RECT 355.705 1.490 355.935 3.325 ;
        RECT 357.225 2.920 357.455 4.350 ;
        RECT 357.945 3.785 358.175 4.580 ;
        RECT 356.190 2.690 357.455 2.920 ;
        RECT 357.945 3.325 359.220 3.555 ;
        RECT 357.225 1.260 357.455 2.390 ;
        RECT 357.945 1.490 358.175 3.325 ;
        RECT 359.465 2.920 359.695 4.350 ;
        RECT 360.185 3.785 360.415 4.580 ;
        RECT 358.430 2.690 359.695 2.920 ;
        RECT 360.185 3.325 361.460 3.555 ;
        RECT 359.465 1.260 359.695 2.390 ;
        RECT 360.185 1.490 360.415 3.325 ;
        RECT 361.705 2.920 361.935 4.350 ;
        RECT 362.570 3.695 362.910 4.580 ;
        RECT 363.545 3.785 363.775 4.580 ;
        RECT 363.545 3.325 364.820 3.555 ;
        RECT 360.670 2.690 361.935 2.920 ;
        RECT 361.705 1.260 361.935 2.390 ;
        RECT 362.570 1.260 362.910 2.950 ;
        RECT 363.545 1.490 363.775 3.325 ;
        RECT 365.065 2.920 365.295 4.350 ;
        RECT 365.785 3.785 366.015 4.580 ;
        RECT 364.030 2.690 365.295 2.920 ;
        RECT 365.785 3.325 367.060 3.555 ;
        RECT 365.065 1.260 365.295 2.390 ;
        RECT 365.785 1.490 366.015 3.325 ;
        RECT 367.305 2.920 367.535 4.350 ;
        RECT 368.025 3.785 368.255 4.580 ;
        RECT 366.270 2.690 367.535 2.920 ;
        RECT 368.025 3.325 369.300 3.555 ;
        RECT 367.305 1.260 367.535 2.390 ;
        RECT 368.025 1.490 368.255 3.325 ;
        RECT 369.545 2.920 369.775 4.350 ;
        RECT 370.265 3.785 370.495 4.580 ;
        RECT 368.510 2.690 369.775 2.920 ;
        RECT 370.265 3.325 371.540 3.555 ;
        RECT 369.545 1.260 369.775 2.390 ;
        RECT 370.265 1.490 370.495 3.325 ;
        RECT 371.785 2.920 372.015 4.350 ;
        RECT 372.505 3.785 372.735 4.580 ;
        RECT 370.750 2.690 372.015 2.920 ;
        RECT 372.505 3.325 373.780 3.555 ;
        RECT 371.785 1.260 372.015 2.390 ;
        RECT 372.505 1.490 372.735 3.325 ;
        RECT 374.025 2.920 374.255 4.350 ;
        RECT 374.745 3.785 374.975 4.580 ;
        RECT 372.990 2.690 374.255 2.920 ;
        RECT 374.745 3.325 376.020 3.555 ;
        RECT 374.025 1.260 374.255 2.390 ;
        RECT 374.745 1.490 374.975 3.325 ;
        RECT 376.265 2.920 376.495 4.350 ;
        RECT 376.985 3.785 377.215 4.580 ;
        RECT 375.230 2.690 376.495 2.920 ;
        RECT 376.985 3.325 378.260 3.555 ;
        RECT 376.265 1.260 376.495 2.390 ;
        RECT 376.985 1.490 377.215 3.325 ;
        RECT 378.505 2.920 378.735 4.350 ;
        RECT 379.225 3.785 379.455 4.580 ;
        RECT 377.470 2.690 378.735 2.920 ;
        RECT 379.225 3.325 380.500 3.555 ;
        RECT 378.505 1.260 378.735 2.390 ;
        RECT 379.225 1.490 379.455 3.325 ;
        RECT 380.745 2.920 380.975 4.350 ;
        RECT 381.465 3.785 381.695 4.580 ;
        RECT 379.710 2.690 380.975 2.920 ;
        RECT 381.465 3.325 382.740 3.555 ;
        RECT 380.745 1.260 380.975 2.390 ;
        RECT 381.465 1.490 381.695 3.325 ;
        RECT 382.985 2.920 383.215 4.350 ;
        RECT 383.850 3.695 384.190 4.580 ;
        RECT 384.825 3.785 385.055 4.580 ;
        RECT 384.825 3.325 386.100 3.555 ;
        RECT 381.950 2.690 383.215 2.920 ;
        RECT 382.985 1.260 383.215 2.390 ;
        RECT 383.850 1.260 384.190 2.950 ;
        RECT 384.825 1.490 385.055 3.325 ;
        RECT 386.345 2.920 386.575 4.350 ;
        RECT 387.065 3.785 387.295 4.580 ;
        RECT 385.310 2.690 386.575 2.920 ;
        RECT 387.065 3.325 388.340 3.555 ;
        RECT 386.345 1.260 386.575 2.390 ;
        RECT 387.065 1.490 387.295 3.325 ;
        RECT 388.585 2.920 388.815 4.350 ;
        RECT 389.305 3.785 389.535 4.580 ;
        RECT 387.550 2.690 388.815 2.920 ;
        RECT 389.305 3.325 390.580 3.555 ;
        RECT 388.585 1.260 388.815 2.390 ;
        RECT 389.305 1.490 389.535 3.325 ;
        RECT 390.825 2.920 391.055 4.350 ;
        RECT 391.545 3.785 391.775 4.580 ;
        RECT 389.790 2.690 391.055 2.920 ;
        RECT 391.545 3.325 392.820 3.555 ;
        RECT 390.825 1.260 391.055 2.390 ;
        RECT 391.545 1.490 391.775 3.325 ;
        RECT 393.065 2.920 393.295 4.350 ;
        RECT 393.785 3.785 394.015 4.580 ;
        RECT 392.030 2.690 393.295 2.920 ;
        RECT 393.785 3.325 395.060 3.555 ;
        RECT 393.065 1.260 393.295 2.390 ;
        RECT 393.785 1.490 394.015 3.325 ;
        RECT 395.305 2.920 395.535 4.350 ;
        RECT 394.270 2.690 395.535 2.920 ;
        RECT 395.305 1.260 395.535 2.390 ;
        RECT 396.025 2.300 396.255 4.080 ;
        RECT 396.485 3.250 397.000 4.230 ;
        RECT 397.365 4.015 397.595 4.580 ;
        RECT 398.110 3.280 398.735 4.305 ;
        RECT 399.385 3.785 399.615 4.580 ;
        RECT 396.485 2.690 397.370 3.250 ;
        RECT 397.750 2.300 398.035 3.050 ;
        RECT 396.025 2.065 398.035 2.300 ;
        RECT 396.025 1.490 396.410 2.065 ;
        RECT 397.310 1.260 397.650 1.750 ;
        RECT 398.265 1.500 398.735 3.280 ;
        RECT 399.385 3.325 400.660 3.555 ;
        RECT 399.385 1.490 399.615 3.325 ;
        RECT 400.905 2.920 401.135 4.350 ;
        RECT 401.625 3.785 401.855 4.580 ;
        RECT 399.870 2.690 401.135 2.920 ;
        RECT 401.625 3.325 402.900 3.555 ;
        RECT 400.905 1.260 401.135 2.390 ;
        RECT 401.625 1.490 401.855 3.325 ;
        RECT 403.145 2.920 403.375 4.350 ;
        RECT 404.010 3.695 404.350 4.580 ;
        RECT 404.985 3.785 405.215 4.580 ;
        RECT 404.985 3.325 406.260 3.555 ;
        RECT 402.110 2.690 403.375 2.920 ;
        RECT 403.145 1.260 403.375 2.390 ;
        RECT 404.010 1.260 404.350 2.950 ;
        RECT 404.985 1.490 405.215 3.325 ;
        RECT 406.505 2.920 406.735 4.350 ;
        RECT 407.225 3.785 407.455 4.580 ;
        RECT 405.470 2.690 406.735 2.920 ;
        RECT 407.225 3.325 408.500 3.555 ;
        RECT 406.505 1.260 406.735 2.390 ;
        RECT 407.225 1.490 407.455 3.325 ;
        RECT 408.745 2.920 408.975 4.350 ;
        RECT 409.465 3.785 409.695 4.580 ;
        RECT 407.710 2.690 408.975 2.920 ;
        RECT 409.465 3.325 410.740 3.555 ;
        RECT 408.745 1.260 408.975 2.390 ;
        RECT 409.465 1.490 409.695 3.325 ;
        RECT 410.985 2.920 411.215 4.350 ;
        RECT 411.705 3.785 411.935 4.580 ;
        RECT 409.950 2.690 411.215 2.920 ;
        RECT 411.705 3.325 412.980 3.555 ;
        RECT 410.985 1.260 411.215 2.390 ;
        RECT 411.705 1.490 411.935 3.325 ;
        RECT 413.225 2.920 413.455 4.350 ;
        RECT 413.945 3.785 414.175 4.580 ;
        RECT 412.190 2.690 413.455 2.920 ;
        RECT 413.945 3.325 415.220 3.555 ;
        RECT 413.225 1.260 413.455 2.390 ;
        RECT 413.945 1.490 414.175 3.325 ;
        RECT 415.465 2.920 415.695 4.350 ;
        RECT 416.185 3.785 416.415 4.580 ;
        RECT 414.430 2.690 415.695 2.920 ;
        RECT 416.185 3.325 417.460 3.555 ;
        RECT 415.465 1.260 415.695 2.390 ;
        RECT 416.185 1.490 416.415 3.325 ;
        RECT 417.705 2.920 417.935 4.350 ;
        RECT 418.425 3.785 418.655 4.580 ;
        RECT 416.670 2.690 417.935 2.920 ;
        RECT 418.425 3.325 419.700 3.555 ;
        RECT 417.705 1.260 417.935 2.390 ;
        RECT 418.425 1.490 418.655 3.325 ;
        RECT 419.945 2.920 420.175 4.350 ;
        RECT 420.665 3.785 420.895 4.580 ;
        RECT 418.910 2.690 420.175 2.920 ;
        RECT 420.665 3.325 421.940 3.555 ;
        RECT 419.945 1.260 420.175 2.390 ;
        RECT 420.665 1.490 420.895 3.325 ;
        RECT 422.185 2.920 422.415 4.350 ;
        RECT 422.905 3.785 423.135 4.580 ;
        RECT 421.150 2.690 422.415 2.920 ;
        RECT 422.905 3.325 424.180 3.555 ;
        RECT 422.185 1.260 422.415 2.390 ;
        RECT 422.905 1.490 423.135 3.325 ;
        RECT 424.425 2.920 424.655 4.350 ;
        RECT 425.290 3.695 425.630 4.580 ;
        RECT 426.265 3.785 426.495 4.580 ;
        RECT 426.265 3.325 427.540 3.555 ;
        RECT 423.390 2.690 424.655 2.920 ;
        RECT 424.425 1.260 424.655 2.390 ;
        RECT 425.290 1.260 425.630 2.950 ;
        RECT 426.265 1.490 426.495 3.325 ;
        RECT 427.785 2.920 428.015 4.350 ;
        RECT 428.505 3.785 428.735 4.580 ;
        RECT 426.750 2.690 428.015 2.920 ;
        RECT 428.505 3.325 429.780 3.555 ;
        RECT 427.785 1.260 428.015 2.390 ;
        RECT 428.505 1.490 428.735 3.325 ;
        RECT 430.025 2.920 430.255 4.350 ;
        RECT 430.745 3.785 430.975 4.580 ;
        RECT 428.990 2.690 430.255 2.920 ;
        RECT 430.745 3.325 432.020 3.555 ;
        RECT 430.025 1.260 430.255 2.390 ;
        RECT 430.745 1.490 430.975 3.325 ;
        RECT 432.265 2.920 432.495 4.350 ;
        RECT 432.985 3.785 433.215 4.580 ;
        RECT 431.230 2.690 432.495 2.920 ;
        RECT 432.985 3.325 434.260 3.555 ;
        RECT 432.265 1.260 432.495 2.390 ;
        RECT 432.985 1.490 433.215 3.325 ;
        RECT 434.505 2.920 434.735 4.350 ;
        RECT 435.225 3.785 435.455 4.580 ;
        RECT 433.470 2.690 434.735 2.920 ;
        RECT 435.225 3.325 436.500 3.555 ;
        RECT 434.505 1.260 434.735 2.390 ;
        RECT 435.225 1.490 435.455 3.325 ;
        RECT 436.745 2.920 436.975 4.350 ;
        RECT 435.710 2.690 436.975 2.920 ;
        RECT 436.745 1.260 436.975 2.390 ;
        RECT 437.465 2.300 437.695 4.080 ;
        RECT 437.925 3.250 438.440 4.230 ;
        RECT 438.805 4.015 439.035 4.580 ;
        RECT 439.550 3.280 440.175 4.305 ;
        RECT 440.825 3.785 441.055 4.580 ;
        RECT 437.925 2.690 438.810 3.250 ;
        RECT 439.190 2.300 439.475 3.050 ;
        RECT 437.465 2.065 439.475 2.300 ;
        RECT 437.465 1.490 437.850 2.065 ;
        RECT 438.750 1.260 439.090 1.750 ;
        RECT 439.705 1.500 440.175 3.280 ;
        RECT 440.825 3.325 442.100 3.555 ;
        RECT 440.825 1.490 441.055 3.325 ;
        RECT 442.345 2.920 442.575 4.350 ;
        RECT 443.065 3.785 443.295 4.580 ;
        RECT 441.310 2.690 442.575 2.920 ;
        RECT 443.065 3.325 444.340 3.555 ;
        RECT 442.345 1.260 442.575 2.390 ;
        RECT 443.065 1.490 443.295 3.325 ;
        RECT 444.585 2.920 444.815 4.350 ;
        RECT 445.450 3.695 445.790 4.580 ;
        RECT 446.425 3.785 446.655 4.580 ;
        RECT 446.425 3.325 447.700 3.555 ;
        RECT 443.550 2.690 444.815 2.920 ;
        RECT 444.585 1.260 444.815 2.390 ;
        RECT 445.450 1.260 445.790 2.950 ;
        RECT 446.425 1.490 446.655 3.325 ;
        RECT 447.945 2.920 448.175 4.350 ;
        RECT 448.665 3.785 448.895 4.580 ;
        RECT 446.910 2.690 448.175 2.920 ;
        RECT 448.665 3.325 449.940 3.555 ;
        RECT 447.945 1.260 448.175 2.390 ;
        RECT 448.665 1.490 448.895 3.325 ;
        RECT 450.185 2.920 450.415 4.350 ;
        RECT 450.905 3.785 451.135 4.580 ;
        RECT 449.150 2.690 450.415 2.920 ;
        RECT 450.905 3.325 452.180 3.555 ;
        RECT 450.185 1.260 450.415 2.390 ;
        RECT 450.905 1.490 451.135 3.325 ;
        RECT 452.425 2.920 452.655 4.350 ;
        RECT 453.145 3.785 453.375 4.580 ;
        RECT 451.390 2.690 452.655 2.920 ;
        RECT 453.145 3.325 454.420 3.555 ;
        RECT 452.425 1.260 452.655 2.390 ;
        RECT 453.145 1.490 453.375 3.325 ;
        RECT 454.665 2.920 454.895 4.350 ;
        RECT 455.385 3.785 455.615 4.580 ;
        RECT 453.630 2.690 454.895 2.920 ;
        RECT 455.385 3.325 456.660 3.555 ;
        RECT 454.665 1.260 454.895 2.390 ;
        RECT 455.385 1.490 455.615 3.325 ;
        RECT 456.905 2.920 457.135 4.350 ;
        RECT 457.625 3.785 457.855 4.580 ;
        RECT 455.870 2.690 457.135 2.920 ;
        RECT 457.625 3.325 458.900 3.555 ;
        RECT 456.905 1.260 457.135 2.390 ;
        RECT 457.625 1.490 457.855 3.325 ;
        RECT 459.145 2.920 459.375 4.350 ;
        RECT 459.865 3.785 460.095 4.580 ;
        RECT 458.110 2.690 459.375 2.920 ;
        RECT 459.865 3.325 461.140 3.555 ;
        RECT 459.145 1.260 459.375 2.390 ;
        RECT 459.865 1.490 460.095 3.325 ;
        RECT 461.385 2.920 461.615 4.350 ;
        RECT 462.105 3.785 462.335 4.580 ;
        RECT 460.350 2.690 461.615 2.920 ;
        RECT 462.105 3.325 463.380 3.555 ;
        RECT 461.385 1.260 461.615 2.390 ;
        RECT 462.105 1.490 462.335 3.325 ;
        RECT 463.625 2.920 463.855 4.350 ;
        RECT 464.345 3.785 464.575 4.580 ;
        RECT 462.590 2.690 463.855 2.920 ;
        RECT 464.345 3.325 465.620 3.555 ;
        RECT 463.625 1.260 463.855 2.390 ;
        RECT 464.345 1.490 464.575 3.325 ;
        RECT 465.865 2.920 466.095 4.350 ;
        RECT 466.730 3.695 467.070 4.580 ;
        RECT 467.705 3.785 467.935 4.580 ;
        RECT 467.705 3.325 468.980 3.555 ;
        RECT 464.830 2.690 466.095 2.920 ;
        RECT 465.865 1.260 466.095 2.390 ;
        RECT 466.730 1.260 467.070 2.950 ;
        RECT 467.705 1.490 467.935 3.325 ;
        RECT 469.225 2.920 469.455 4.350 ;
        RECT 469.945 3.785 470.175 4.580 ;
        RECT 468.190 2.690 469.455 2.920 ;
        RECT 469.945 3.325 471.220 3.555 ;
        RECT 469.225 1.260 469.455 2.390 ;
        RECT 469.945 1.490 470.175 3.325 ;
        RECT 471.465 2.920 471.695 4.350 ;
        RECT 472.185 3.785 472.415 4.580 ;
        RECT 470.430 2.690 471.695 2.920 ;
        RECT 472.185 3.325 473.460 3.555 ;
        RECT 471.465 1.260 471.695 2.390 ;
        RECT 472.185 1.490 472.415 3.325 ;
        RECT 473.705 2.920 473.935 4.350 ;
        RECT 474.425 3.785 474.655 4.580 ;
        RECT 472.670 2.690 473.935 2.920 ;
        RECT 474.425 3.325 475.700 3.555 ;
        RECT 473.705 1.260 473.935 2.390 ;
        RECT 474.425 1.490 474.655 3.325 ;
        RECT 475.945 2.920 476.175 4.350 ;
        RECT 476.665 3.785 476.895 4.580 ;
        RECT 474.910 2.690 476.175 2.920 ;
        RECT 476.665 3.325 477.940 3.555 ;
        RECT 475.945 1.260 476.175 2.390 ;
        RECT 476.665 1.490 476.895 3.325 ;
        RECT 478.185 2.920 478.415 4.350 ;
        RECT 478.905 3.785 479.135 4.580 ;
        RECT 477.150 2.690 478.415 2.920 ;
        RECT 478.905 3.325 480.180 3.555 ;
        RECT 478.185 1.260 478.415 2.390 ;
        RECT 478.905 1.490 479.135 3.325 ;
        RECT 480.425 2.920 480.655 4.350 ;
        RECT 479.390 2.690 480.655 2.920 ;
        RECT 480.425 1.260 480.655 2.390 ;
        RECT 481.145 2.300 481.375 4.080 ;
        RECT 481.605 3.250 482.120 4.230 ;
        RECT 482.485 4.015 482.715 4.580 ;
        RECT 483.230 3.280 483.855 4.305 ;
        RECT 484.505 3.785 484.735 4.580 ;
        RECT 481.605 2.690 482.490 3.250 ;
        RECT 482.870 2.300 483.155 3.050 ;
        RECT 481.145 2.065 483.155 2.300 ;
        RECT 481.145 1.490 481.530 2.065 ;
        RECT 482.430 1.260 482.770 1.750 ;
        RECT 483.385 1.500 483.855 3.280 ;
        RECT 484.505 3.325 485.780 3.555 ;
        RECT 484.505 1.490 484.735 3.325 ;
        RECT 486.025 2.920 486.255 4.350 ;
        RECT 486.890 3.695 487.230 4.580 ;
        RECT 487.865 3.785 488.095 4.580 ;
        RECT 487.865 3.325 489.140 3.555 ;
        RECT 484.990 2.690 486.255 2.920 ;
        RECT 486.025 1.260 486.255 2.390 ;
        RECT 486.890 1.260 487.230 2.950 ;
        RECT 487.865 1.490 488.095 3.325 ;
        RECT 489.385 2.920 489.615 4.350 ;
        RECT 490.105 3.785 490.335 4.580 ;
        RECT 488.350 2.690 489.615 2.920 ;
        RECT 490.105 3.325 491.380 3.555 ;
        RECT 489.385 1.260 489.615 2.390 ;
        RECT 490.105 1.490 490.335 3.325 ;
        RECT 491.625 2.920 491.855 4.350 ;
        RECT 492.345 3.785 492.575 4.580 ;
        RECT 490.590 2.690 491.855 2.920 ;
        RECT 492.345 3.325 493.620 3.555 ;
        RECT 491.625 1.260 491.855 2.390 ;
        RECT 492.345 1.490 492.575 3.325 ;
        RECT 493.865 2.920 494.095 4.350 ;
        RECT 494.585 3.785 494.815 4.580 ;
        RECT 492.830 2.690 494.095 2.920 ;
        RECT 494.585 3.325 495.860 3.555 ;
        RECT 493.865 1.260 494.095 2.390 ;
        RECT 494.585 1.490 494.815 3.325 ;
        RECT 496.105 2.920 496.335 4.350 ;
        RECT 496.825 3.785 497.055 4.580 ;
        RECT 495.070 2.690 496.335 2.920 ;
        RECT 496.825 3.325 498.100 3.555 ;
        RECT 496.105 1.260 496.335 2.390 ;
        RECT 496.825 1.490 497.055 3.325 ;
        RECT 498.345 2.920 498.575 4.350 ;
        RECT 499.065 3.785 499.295 4.580 ;
        RECT 497.310 2.690 498.575 2.920 ;
        RECT 499.065 3.325 500.340 3.555 ;
        RECT 498.345 1.260 498.575 2.390 ;
        RECT 499.065 1.490 499.295 3.325 ;
        RECT 500.585 2.920 500.815 4.350 ;
        RECT 501.305 3.785 501.535 4.580 ;
        RECT 499.550 2.690 500.815 2.920 ;
        RECT 501.305 3.325 502.580 3.555 ;
        RECT 500.585 1.260 500.815 2.390 ;
        RECT 501.305 1.490 501.535 3.325 ;
        RECT 502.825 2.920 503.055 4.350 ;
        RECT 503.545 3.785 503.775 4.580 ;
        RECT 501.790 2.690 503.055 2.920 ;
        RECT 503.545 3.325 504.820 3.555 ;
        RECT 502.825 1.260 503.055 2.390 ;
        RECT 503.545 1.490 503.775 3.325 ;
        RECT 505.065 2.920 505.295 4.350 ;
        RECT 505.785 3.785 506.015 4.580 ;
        RECT 504.030 2.690 505.295 2.920 ;
        RECT 505.785 3.325 507.060 3.555 ;
        RECT 505.065 1.260 505.295 2.390 ;
        RECT 505.785 1.490 506.015 3.325 ;
        RECT 507.305 2.920 507.535 4.350 ;
        RECT 508.170 3.695 508.510 4.580 ;
        RECT 509.145 3.785 509.375 4.580 ;
        RECT 509.145 3.325 510.420 3.555 ;
        RECT 506.270 2.690 507.535 2.920 ;
        RECT 507.305 1.260 507.535 2.390 ;
        RECT 508.170 1.260 508.510 2.950 ;
        RECT 509.145 1.490 509.375 3.325 ;
        RECT 510.665 2.920 510.895 4.350 ;
        RECT 511.385 3.785 511.615 4.580 ;
        RECT 509.630 2.690 510.895 2.920 ;
        RECT 511.385 3.325 512.660 3.555 ;
        RECT 510.665 1.260 510.895 2.390 ;
        RECT 511.385 1.490 511.615 3.325 ;
        RECT 512.905 2.920 513.135 4.350 ;
        RECT 513.625 3.785 513.855 4.580 ;
        RECT 511.870 2.690 513.135 2.920 ;
        RECT 513.625 3.325 514.900 3.555 ;
        RECT 512.905 1.260 513.135 2.390 ;
        RECT 513.625 1.490 513.855 3.325 ;
        RECT 515.145 2.920 515.375 4.350 ;
        RECT 515.865 3.785 516.095 4.580 ;
        RECT 514.110 2.690 515.375 2.920 ;
        RECT 515.865 3.325 517.140 3.555 ;
        RECT 515.145 1.260 515.375 2.390 ;
        RECT 515.865 1.490 516.095 3.325 ;
        RECT 517.385 2.920 517.615 4.350 ;
        RECT 518.105 3.785 518.335 4.580 ;
        RECT 516.350 2.690 517.615 2.920 ;
        RECT 518.105 3.325 519.380 3.555 ;
        RECT 517.385 1.260 517.615 2.390 ;
        RECT 518.105 1.490 518.335 3.325 ;
        RECT 519.625 2.920 519.855 4.350 ;
        RECT 520.345 3.785 520.575 4.580 ;
        RECT 518.590 2.690 519.855 2.920 ;
        RECT 520.345 3.325 521.620 3.555 ;
        RECT 519.625 1.260 519.855 2.390 ;
        RECT 520.345 1.490 520.575 3.325 ;
        RECT 521.865 2.920 522.095 4.350 ;
        RECT 520.830 2.690 522.095 2.920 ;
        RECT 521.865 1.260 522.095 2.390 ;
        RECT 522.585 2.300 522.815 4.080 ;
        RECT 523.045 3.250 523.560 4.230 ;
        RECT 523.925 4.015 524.155 4.580 ;
        RECT 524.670 3.280 525.295 4.305 ;
        RECT 525.945 3.785 526.175 4.580 ;
        RECT 523.045 2.690 523.930 3.250 ;
        RECT 524.310 2.300 524.595 3.050 ;
        RECT 522.585 2.065 524.595 2.300 ;
        RECT 522.585 1.490 522.970 2.065 ;
        RECT 523.870 1.260 524.210 1.750 ;
        RECT 524.825 1.500 525.295 3.280 ;
        RECT 525.945 3.325 527.220 3.555 ;
        RECT 525.945 1.490 526.175 3.325 ;
        RECT 527.465 2.920 527.695 4.350 ;
        RECT 528.330 3.695 528.670 4.580 ;
        RECT 529.305 3.785 529.535 4.580 ;
        RECT 529.305 3.325 530.580 3.555 ;
        RECT 526.430 2.690 527.695 2.920 ;
        RECT 527.465 1.260 527.695 2.390 ;
        RECT 528.330 1.260 528.670 2.950 ;
        RECT 529.305 1.490 529.535 3.325 ;
        RECT 530.825 2.920 531.055 4.350 ;
        RECT 531.545 3.785 531.775 4.580 ;
        RECT 529.790 2.690 531.055 2.920 ;
        RECT 531.545 3.325 532.820 3.555 ;
        RECT 530.825 1.260 531.055 2.390 ;
        RECT 531.545 1.490 531.775 3.325 ;
        RECT 533.065 2.920 533.295 4.350 ;
        RECT 533.785 3.785 534.015 4.580 ;
        RECT 532.030 2.690 533.295 2.920 ;
        RECT 533.785 3.325 535.060 3.555 ;
        RECT 533.065 1.260 533.295 2.390 ;
        RECT 533.785 1.490 534.015 3.325 ;
        RECT 535.305 2.920 535.535 4.350 ;
        RECT 536.025 3.785 536.255 4.580 ;
        RECT 534.270 2.690 535.535 2.920 ;
        RECT 536.025 3.325 537.300 3.555 ;
        RECT 535.305 1.260 535.535 2.390 ;
        RECT 536.025 1.490 536.255 3.325 ;
        RECT 537.545 2.920 537.775 4.350 ;
        RECT 538.265 3.785 538.495 4.580 ;
        RECT 536.510 2.690 537.775 2.920 ;
        RECT 538.265 3.325 539.540 3.555 ;
        RECT 537.545 1.260 537.775 2.390 ;
        RECT 538.265 1.490 538.495 3.325 ;
        RECT 539.785 2.920 540.015 4.350 ;
        RECT 540.505 3.785 540.735 4.580 ;
        RECT 538.750 2.690 540.015 2.920 ;
        RECT 540.505 3.325 541.780 3.555 ;
        RECT 539.785 1.260 540.015 2.390 ;
        RECT 540.505 1.490 540.735 3.325 ;
        RECT 542.025 2.920 542.255 4.350 ;
        RECT 542.745 3.785 542.975 4.580 ;
        RECT 540.990 2.690 542.255 2.920 ;
        RECT 542.745 3.325 544.020 3.555 ;
        RECT 542.025 1.260 542.255 2.390 ;
        RECT 542.745 1.490 542.975 3.325 ;
        RECT 544.265 2.920 544.495 4.350 ;
        RECT 544.985 3.785 545.215 4.580 ;
        RECT 543.230 2.690 544.495 2.920 ;
        RECT 544.985 3.325 546.260 3.555 ;
        RECT 544.265 1.260 544.495 2.390 ;
        RECT 544.985 1.490 545.215 3.325 ;
        RECT 546.505 2.920 546.735 4.350 ;
        RECT 547.225 3.785 547.455 4.580 ;
        RECT 545.470 2.690 546.735 2.920 ;
        RECT 547.225 3.325 548.500 3.555 ;
        RECT 546.505 1.260 546.735 2.390 ;
        RECT 547.225 1.490 547.455 3.325 ;
        RECT 548.745 2.920 548.975 4.350 ;
        RECT 549.610 3.695 549.950 4.580 ;
        RECT 550.585 3.785 550.815 4.580 ;
        RECT 550.585 3.325 551.860 3.555 ;
        RECT 547.710 2.690 548.975 2.920 ;
        RECT 548.745 1.260 548.975 2.390 ;
        RECT 549.610 1.260 549.950 2.950 ;
        RECT 550.585 1.490 550.815 3.325 ;
        RECT 552.105 2.920 552.335 4.350 ;
        RECT 552.825 3.785 553.055 4.580 ;
        RECT 551.070 2.690 552.335 2.920 ;
        RECT 552.825 3.325 554.100 3.555 ;
        RECT 552.105 1.260 552.335 2.390 ;
        RECT 552.825 1.490 553.055 3.325 ;
        RECT 554.345 2.920 554.575 4.350 ;
        RECT 555.065 3.785 555.295 4.580 ;
        RECT 553.310 2.690 554.575 2.920 ;
        RECT 555.065 3.325 556.340 3.555 ;
        RECT 554.345 1.260 554.575 2.390 ;
        RECT 555.065 1.490 555.295 3.325 ;
        RECT 556.585 2.920 556.815 4.350 ;
        RECT 557.305 3.785 557.535 4.580 ;
        RECT 555.550 2.690 556.815 2.920 ;
        RECT 557.305 3.325 558.580 3.555 ;
        RECT 556.585 1.260 556.815 2.390 ;
        RECT 557.305 1.490 557.535 3.325 ;
        RECT 558.825 2.920 559.055 4.350 ;
        RECT 559.545 3.785 559.775 4.580 ;
        RECT 557.790 2.690 559.055 2.920 ;
        RECT 559.545 3.325 560.820 3.555 ;
        RECT 558.825 1.260 559.055 2.390 ;
        RECT 559.545 1.490 559.775 3.325 ;
        RECT 561.065 2.920 561.295 4.350 ;
        RECT 561.785 3.785 562.015 4.580 ;
        RECT 560.030 2.690 561.295 2.920 ;
        RECT 561.785 3.325 563.060 3.555 ;
        RECT 561.065 1.260 561.295 2.390 ;
        RECT 561.785 1.490 562.015 3.325 ;
        RECT 563.305 2.920 563.535 4.350 ;
        RECT 564.025 3.785 564.255 4.580 ;
        RECT 562.270 2.690 563.535 2.920 ;
        RECT 564.025 3.325 565.300 3.555 ;
        RECT 563.305 1.260 563.535 2.390 ;
        RECT 564.025 1.490 564.255 3.325 ;
        RECT 565.545 2.920 565.775 4.350 ;
        RECT 564.510 2.690 565.775 2.920 ;
        RECT 565.545 1.260 565.775 2.390 ;
        RECT 566.265 2.300 566.495 4.080 ;
        RECT 566.725 3.250 567.240 4.230 ;
        RECT 567.605 4.015 567.835 4.580 ;
        RECT 568.350 3.280 568.975 4.305 ;
        RECT 569.770 3.695 570.110 4.580 ;
        RECT 570.745 3.785 570.975 4.580 ;
        RECT 566.725 2.690 567.610 3.250 ;
        RECT 567.990 2.300 568.275 3.050 ;
        RECT 566.265 2.065 568.275 2.300 ;
        RECT 566.265 1.490 566.650 2.065 ;
        RECT 567.550 1.260 567.890 1.750 ;
        RECT 568.505 1.500 568.975 3.280 ;
        RECT 570.745 3.325 572.020 3.555 ;
        RECT 569.770 1.260 570.110 2.950 ;
        RECT 570.745 1.490 570.975 3.325 ;
        RECT 572.265 2.920 572.495 4.350 ;
        RECT 572.985 3.785 573.215 4.580 ;
        RECT 571.230 2.690 572.495 2.920 ;
        RECT 572.985 3.325 574.260 3.555 ;
        RECT 572.265 1.260 572.495 2.390 ;
        RECT 572.985 1.490 573.215 3.325 ;
        RECT 574.505 2.920 574.735 4.350 ;
        RECT 575.225 3.785 575.455 4.580 ;
        RECT 573.470 2.690 574.735 2.920 ;
        RECT 575.225 3.325 576.500 3.555 ;
        RECT 574.505 1.260 574.735 2.390 ;
        RECT 575.225 1.490 575.455 3.325 ;
        RECT 576.745 2.920 576.975 4.350 ;
        RECT 577.465 3.785 577.695 4.580 ;
        RECT 575.710 2.690 576.975 2.920 ;
        RECT 577.465 3.325 578.740 3.555 ;
        RECT 576.745 1.260 576.975 2.390 ;
        RECT 577.465 1.490 577.695 3.325 ;
        RECT 578.985 2.920 579.215 4.350 ;
        RECT 579.705 3.785 579.935 4.580 ;
        RECT 577.950 2.690 579.215 2.920 ;
        RECT 579.705 3.325 580.980 3.555 ;
        RECT 578.985 1.260 579.215 2.390 ;
        RECT 579.705 1.490 579.935 3.325 ;
        RECT 581.225 2.920 581.455 4.350 ;
        RECT 581.945 3.785 582.175 4.580 ;
        RECT 580.190 2.690 581.455 2.920 ;
        RECT 581.945 3.325 583.220 3.555 ;
        RECT 581.225 1.260 581.455 2.390 ;
        RECT 581.945 1.490 582.175 3.325 ;
        RECT 583.465 2.920 583.695 4.350 ;
        RECT 584.185 3.785 584.415 4.580 ;
        RECT 582.430 2.690 583.695 2.920 ;
        RECT 584.185 3.325 585.460 3.555 ;
        RECT 583.465 1.260 583.695 2.390 ;
        RECT 584.185 1.490 584.415 3.325 ;
        RECT 585.705 2.920 585.935 4.350 ;
        RECT 586.425 3.785 586.655 4.580 ;
        RECT 584.670 2.690 585.935 2.920 ;
        RECT 586.425 3.325 587.700 3.555 ;
        RECT 585.705 1.260 585.935 2.390 ;
        RECT 586.425 1.490 586.655 3.325 ;
        RECT 587.945 2.920 588.175 4.350 ;
        RECT 588.665 3.785 588.895 4.580 ;
        RECT 586.910 2.690 588.175 2.920 ;
        RECT 588.665 3.325 589.940 3.555 ;
        RECT 587.945 1.260 588.175 2.390 ;
        RECT 588.665 1.490 588.895 3.325 ;
        RECT 590.185 2.920 590.415 4.350 ;
        RECT 591.050 3.695 591.390 4.580 ;
        RECT 592.025 3.785 592.255 4.580 ;
        RECT 592.025 3.325 593.300 3.555 ;
        RECT 589.150 2.690 590.415 2.920 ;
        RECT 590.185 1.260 590.415 2.390 ;
        RECT 591.050 1.260 591.390 2.950 ;
        RECT 592.025 1.490 592.255 3.325 ;
        RECT 593.545 2.920 593.775 4.350 ;
        RECT 594.265 3.785 594.495 4.580 ;
        RECT 592.510 2.690 593.775 2.920 ;
        RECT 594.265 3.325 595.540 3.555 ;
        RECT 593.545 1.260 593.775 2.390 ;
        RECT 594.265 1.490 594.495 3.325 ;
        RECT 595.785 2.920 596.015 4.350 ;
        RECT 596.505 3.785 596.735 4.580 ;
        RECT 594.750 2.690 596.015 2.920 ;
        RECT 596.505 3.325 597.780 3.555 ;
        RECT 595.785 1.260 596.015 2.390 ;
        RECT 596.505 1.490 596.735 3.325 ;
        RECT 598.025 2.920 598.255 4.350 ;
        RECT 598.745 3.785 598.975 4.580 ;
        RECT 596.990 2.690 598.255 2.920 ;
        RECT 598.745 3.325 600.020 3.555 ;
        RECT 598.025 1.260 598.255 2.390 ;
        RECT 598.745 1.490 598.975 3.325 ;
        RECT 600.265 2.920 600.495 4.350 ;
        RECT 600.985 3.785 601.215 4.580 ;
        RECT 599.230 2.690 600.495 2.920 ;
        RECT 600.985 3.325 602.260 3.555 ;
        RECT 600.265 1.260 600.495 2.390 ;
        RECT 600.985 1.490 601.215 3.325 ;
        RECT 602.505 2.920 602.735 4.350 ;
        RECT 603.225 3.785 603.455 4.580 ;
        RECT 601.470 2.690 602.735 2.920 ;
        RECT 603.225 3.325 604.500 3.555 ;
        RECT 602.505 1.260 602.735 2.390 ;
        RECT 603.225 1.490 603.455 3.325 ;
        RECT 604.745 2.920 604.975 4.350 ;
        RECT 605.465 3.785 605.695 4.580 ;
        RECT 603.710 2.690 604.975 2.920 ;
        RECT 605.465 3.325 606.740 3.555 ;
        RECT 604.745 1.260 604.975 2.390 ;
        RECT 605.465 1.490 605.695 3.325 ;
        RECT 606.985 2.920 607.215 4.350 ;
        RECT 605.950 2.690 607.215 2.920 ;
        RECT 606.985 1.260 607.215 2.390 ;
        RECT 607.705 2.300 607.935 4.080 ;
        RECT 608.165 3.250 608.680 4.230 ;
        RECT 609.045 4.015 609.275 4.580 ;
        RECT 609.790 3.280 610.415 4.305 ;
        RECT 611.210 3.695 611.550 4.580 ;
        RECT 612.185 3.785 612.415 4.580 ;
        RECT 608.165 2.690 609.050 3.250 ;
        RECT 609.430 2.300 609.715 3.050 ;
        RECT 607.705 2.065 609.715 2.300 ;
        RECT 607.705 1.490 608.090 2.065 ;
        RECT 608.990 1.260 609.330 1.750 ;
        RECT 609.945 1.500 610.415 3.280 ;
        RECT 612.185 3.325 613.460 3.555 ;
        RECT 611.210 1.260 611.550 2.950 ;
        RECT 612.185 1.490 612.415 3.325 ;
        RECT 613.705 2.920 613.935 4.350 ;
        RECT 614.425 3.785 614.655 4.580 ;
        RECT 612.670 2.690 613.935 2.920 ;
        RECT 614.425 3.325 615.700 3.555 ;
        RECT 613.705 1.260 613.935 2.390 ;
        RECT 614.425 1.490 614.655 3.325 ;
        RECT 615.945 2.920 616.175 4.350 ;
        RECT 616.665 3.785 616.895 4.580 ;
        RECT 614.910 2.690 616.175 2.920 ;
        RECT 616.665 3.325 617.940 3.555 ;
        RECT 615.945 1.260 616.175 2.390 ;
        RECT 616.665 1.490 616.895 3.325 ;
        RECT 618.185 2.920 618.415 4.350 ;
        RECT 618.905 3.785 619.135 4.580 ;
        RECT 617.150 2.690 618.415 2.920 ;
        RECT 618.905 3.325 620.180 3.555 ;
        RECT 618.185 1.260 618.415 2.390 ;
        RECT 618.905 1.490 619.135 3.325 ;
        RECT 620.425 2.920 620.655 4.350 ;
        RECT 621.145 3.785 621.375 4.580 ;
        RECT 619.390 2.690 620.655 2.920 ;
        RECT 621.145 3.325 622.420 3.555 ;
        RECT 620.425 1.260 620.655 2.390 ;
        RECT 621.145 1.490 621.375 3.325 ;
        RECT 622.665 2.920 622.895 4.350 ;
        RECT 623.385 3.785 623.615 4.580 ;
        RECT 621.630 2.690 622.895 2.920 ;
        RECT 623.385 3.325 624.660 3.555 ;
        RECT 622.665 1.260 622.895 2.390 ;
        RECT 623.385 1.490 623.615 3.325 ;
        RECT 624.905 2.920 625.135 4.350 ;
        RECT 625.625 3.785 625.855 4.580 ;
        RECT 623.870 2.690 625.135 2.920 ;
        RECT 625.625 3.325 626.900 3.555 ;
        RECT 624.905 1.260 625.135 2.390 ;
        RECT 625.625 1.490 625.855 3.325 ;
        RECT 627.145 2.920 627.375 4.350 ;
        RECT 627.865 3.785 628.095 4.580 ;
        RECT 626.110 2.690 627.375 2.920 ;
        RECT 627.865 3.325 629.140 3.555 ;
        RECT 627.145 1.260 627.375 2.390 ;
        RECT 627.865 1.490 628.095 3.325 ;
        RECT 629.385 2.920 629.615 4.350 ;
        RECT 630.105 3.785 630.335 4.580 ;
        RECT 628.350 2.690 629.615 2.920 ;
        RECT 630.105 3.325 631.380 3.555 ;
        RECT 629.385 1.260 629.615 2.390 ;
        RECT 630.105 1.490 630.335 3.325 ;
        RECT 631.625 2.920 631.855 4.350 ;
        RECT 632.490 3.695 632.830 4.580 ;
        RECT 633.465 3.785 633.695 4.580 ;
        RECT 633.465 3.325 634.740 3.555 ;
        RECT 630.590 2.690 631.855 2.920 ;
        RECT 631.625 1.260 631.855 2.390 ;
        RECT 632.490 1.260 632.830 2.950 ;
        RECT 633.465 1.490 633.695 3.325 ;
        RECT 634.985 2.920 635.215 4.350 ;
        RECT 635.705 3.785 635.935 4.580 ;
        RECT 633.950 2.690 635.215 2.920 ;
        RECT 635.705 3.325 636.980 3.555 ;
        RECT 634.985 1.260 635.215 2.390 ;
        RECT 635.705 1.490 635.935 3.325 ;
        RECT 637.225 2.920 637.455 4.350 ;
        RECT 637.945 3.785 638.175 4.580 ;
        RECT 636.190 2.690 637.455 2.920 ;
        RECT 637.945 3.325 639.220 3.555 ;
        RECT 637.225 1.260 637.455 2.390 ;
        RECT 637.945 1.490 638.175 3.325 ;
        RECT 639.465 2.920 639.695 4.350 ;
        RECT 640.185 3.785 640.415 4.580 ;
        RECT 638.430 2.690 639.695 2.920 ;
        RECT 640.185 3.325 641.460 3.555 ;
        RECT 639.465 1.260 639.695 2.390 ;
        RECT 640.185 1.490 640.415 3.325 ;
        RECT 641.705 2.920 641.935 4.350 ;
        RECT 642.425 3.785 642.655 4.580 ;
        RECT 640.670 2.690 641.935 2.920 ;
        RECT 642.425 3.325 643.700 3.555 ;
        RECT 641.705 1.260 641.935 2.390 ;
        RECT 642.425 1.490 642.655 3.325 ;
        RECT 643.945 2.920 644.175 4.350 ;
        RECT 644.665 3.785 644.895 4.580 ;
        RECT 642.910 2.690 644.175 2.920 ;
        RECT 644.665 3.325 645.940 3.555 ;
        RECT 643.945 1.260 644.175 2.390 ;
        RECT 644.665 1.490 644.895 3.325 ;
        RECT 646.185 2.920 646.415 4.350 ;
        RECT 646.905 3.785 647.135 4.580 ;
        RECT 645.150 2.690 646.415 2.920 ;
        RECT 646.905 3.325 648.180 3.555 ;
        RECT 646.185 1.260 646.415 2.390 ;
        RECT 646.905 1.490 647.135 3.325 ;
        RECT 648.425 2.920 648.655 4.350 ;
        RECT 649.145 3.785 649.375 4.580 ;
        RECT 647.390 2.690 648.655 2.920 ;
        RECT 649.145 3.325 650.420 3.555 ;
        RECT 648.425 1.260 648.655 2.390 ;
        RECT 649.145 1.490 649.375 3.325 ;
        RECT 650.665 2.920 650.895 4.350 ;
        RECT 649.630 2.690 650.895 2.920 ;
        RECT 650.665 1.260 650.895 2.390 ;
        RECT 651.385 2.300 651.615 4.080 ;
        RECT 651.845 3.250 652.360 4.230 ;
        RECT 652.725 4.015 652.955 4.580 ;
        RECT 653.470 3.280 654.095 4.305 ;
        RECT 654.890 3.695 655.230 4.580 ;
        RECT 655.865 3.785 656.095 4.580 ;
        RECT 651.845 2.690 652.730 3.250 ;
        RECT 653.110 2.300 653.395 3.050 ;
        RECT 651.385 2.065 653.395 2.300 ;
        RECT 651.385 1.490 651.770 2.065 ;
        RECT 652.670 1.260 653.010 1.750 ;
        RECT 653.625 1.500 654.095 3.280 ;
        RECT 655.865 3.325 657.140 3.555 ;
        RECT 654.890 1.260 655.230 2.950 ;
        RECT 655.865 1.490 656.095 3.325 ;
        RECT 657.385 2.920 657.615 4.350 ;
        RECT 658.105 3.785 658.335 4.580 ;
        RECT 656.350 2.690 657.615 2.920 ;
        RECT 658.105 3.325 659.380 3.555 ;
        RECT 657.385 1.260 657.615 2.390 ;
        RECT 658.105 1.490 658.335 3.325 ;
        RECT 659.625 2.920 659.855 4.350 ;
        RECT 660.345 3.785 660.575 4.580 ;
        RECT 658.590 2.690 659.855 2.920 ;
        RECT 660.345 3.325 661.620 3.555 ;
        RECT 659.625 1.260 659.855 2.390 ;
        RECT 660.345 1.490 660.575 3.325 ;
        RECT 661.865 2.920 662.095 4.350 ;
        RECT 662.585 3.785 662.815 4.580 ;
        RECT 660.830 2.690 662.095 2.920 ;
        RECT 662.585 3.325 663.860 3.555 ;
        RECT 661.865 1.260 662.095 2.390 ;
        RECT 662.585 1.490 662.815 3.325 ;
        RECT 664.105 2.920 664.335 4.350 ;
        RECT 664.825 3.785 665.055 4.580 ;
        RECT 663.070 2.690 664.335 2.920 ;
        RECT 664.825 3.325 666.100 3.555 ;
        RECT 664.105 1.260 664.335 2.390 ;
        RECT 664.825 1.490 665.055 3.325 ;
        RECT 666.345 2.920 666.575 4.350 ;
        RECT 667.065 3.785 667.295 4.580 ;
        RECT 665.310 2.690 666.575 2.920 ;
        RECT 667.065 3.325 668.340 3.555 ;
        RECT 666.345 1.260 666.575 2.390 ;
        RECT 667.065 1.490 667.295 3.325 ;
        RECT 668.585 2.920 668.815 4.350 ;
        RECT 669.305 3.785 669.535 4.580 ;
        RECT 667.550 2.690 668.815 2.920 ;
        RECT 669.305 3.325 670.580 3.555 ;
        RECT 668.585 1.260 668.815 2.390 ;
        RECT 669.305 1.490 669.535 3.325 ;
        RECT 670.825 2.920 671.055 4.350 ;
        RECT 671.545 3.785 671.775 4.580 ;
        RECT 669.790 2.690 671.055 2.920 ;
        RECT 671.545 3.325 672.820 3.555 ;
        RECT 670.825 1.260 671.055 2.390 ;
        RECT 671.545 1.490 671.775 3.325 ;
        RECT 673.065 2.920 673.295 4.350 ;
        RECT 673.785 3.785 674.015 4.580 ;
        RECT 672.030 2.690 673.295 2.920 ;
        RECT 673.785 3.325 675.060 3.555 ;
        RECT 673.065 1.260 673.295 2.390 ;
        RECT 673.785 1.490 674.015 3.325 ;
        RECT 675.305 2.920 675.535 4.350 ;
        RECT 676.170 3.695 676.510 4.580 ;
        RECT 677.145 3.785 677.375 4.580 ;
        RECT 677.145 3.325 678.420 3.555 ;
        RECT 674.270 2.690 675.535 2.920 ;
        RECT 675.305 1.260 675.535 2.390 ;
        RECT 676.170 1.260 676.510 2.950 ;
        RECT 677.145 1.490 677.375 3.325 ;
        RECT 678.665 2.920 678.895 4.350 ;
        RECT 679.510 3.690 679.850 4.580 ;
        RECT 677.630 2.690 678.895 2.920 ;
        RECT 678.665 1.260 678.895 2.390 ;
        RECT 679.510 1.260 679.850 2.960 ;
        RECT 122.090 0.660 680.260 1.260 ;
        RECT 122.090 0.610 122.470 0.660 ;
        RECT 122.820 0.620 123.260 0.660 ;
      LAYER Via1 ;
        RECT 2.190 59.990 2.450 60.250 ;
        RECT 20.035 59.990 20.295 60.250 ;
        RECT 0.825 58.805 1.085 59.065 ;
        RECT 0.825 58.145 1.085 58.405 ;
        RECT 0.825 57.485 1.085 57.745 ;
        RECT 0.825 56.825 1.085 57.085 ;
        RECT 0.825 56.165 1.085 56.425 ;
        RECT 0.825 55.505 1.085 55.765 ;
        RECT 0.825 54.845 1.085 55.105 ;
        RECT 0.825 54.185 1.085 54.445 ;
        RECT 0.825 53.525 1.085 53.785 ;
        RECT 0.825 52.865 1.085 53.125 ;
        RECT 0.825 52.205 1.085 52.465 ;
        RECT 0.825 51.545 1.085 51.805 ;
        RECT 0.825 50.885 1.085 51.145 ;
        RECT 0.825 50.225 1.085 50.485 ;
        RECT 5.310 47.865 5.570 48.125 ;
        RECT 5.970 47.865 6.230 48.125 ;
        RECT 6.630 47.865 6.890 48.125 ;
        RECT 5.310 47.205 5.570 47.465 ;
        RECT 5.970 47.205 6.230 47.465 ;
        RECT 6.630 47.205 6.890 47.465 ;
        RECT 5.310 46.545 5.570 46.805 ;
        RECT 5.970 46.545 6.230 46.805 ;
        RECT 6.630 46.545 6.890 46.805 ;
        RECT 5.310 22.265 5.570 22.525 ;
        RECT 5.970 22.265 6.230 22.525 ;
        RECT 6.630 22.265 6.890 22.525 ;
        RECT 5.310 21.605 5.570 21.865 ;
        RECT 5.970 21.605 6.230 21.865 ;
        RECT 6.630 21.605 6.890 21.865 ;
        RECT 5.310 20.945 5.570 21.205 ;
        RECT 5.970 20.945 6.230 21.205 ;
        RECT 6.630 20.945 6.890 21.205 ;
        RECT 11.115 58.805 11.375 59.065 ;
        RECT 11.115 58.145 11.375 58.405 ;
        RECT 11.115 57.485 11.375 57.745 ;
        RECT 11.115 56.825 11.375 57.085 ;
        RECT 11.115 56.165 11.375 56.425 ;
        RECT 11.115 55.505 11.375 55.765 ;
        RECT 11.115 54.845 11.375 55.105 ;
        RECT 11.115 54.185 11.375 54.445 ;
        RECT 11.115 53.525 11.375 53.785 ;
        RECT 11.115 52.865 11.375 53.125 ;
        RECT 11.115 52.205 11.375 52.465 ;
        RECT 11.115 51.545 11.375 51.805 ;
        RECT 11.115 50.885 11.375 51.145 ;
        RECT 11.115 50.225 11.375 50.485 ;
        RECT 22.765 59.990 23.025 60.250 ;
        RECT 40.610 59.990 40.870 60.250 ;
        RECT 15.610 45.165 15.870 45.425 ;
        RECT 16.270 45.165 16.530 45.425 ;
        RECT 16.930 45.165 17.190 45.425 ;
        RECT 15.610 44.505 15.870 44.765 ;
        RECT 16.270 44.505 16.530 44.765 ;
        RECT 16.930 44.505 17.190 44.765 ;
        RECT 15.610 43.845 15.870 44.105 ;
        RECT 16.270 43.845 16.530 44.105 ;
        RECT 16.930 43.845 17.190 44.105 ;
        RECT 15.610 24.965 15.870 25.225 ;
        RECT 16.270 24.965 16.530 25.225 ;
        RECT 16.930 24.965 17.190 25.225 ;
        RECT 15.610 24.305 15.870 24.565 ;
        RECT 16.270 24.305 16.530 24.565 ;
        RECT 16.930 24.305 17.190 24.565 ;
        RECT 15.610 23.645 15.870 23.905 ;
        RECT 16.270 23.645 16.530 23.905 ;
        RECT 16.930 23.645 17.190 23.905 ;
        RECT 9.750 8.805 10.010 9.065 ;
        RECT 21.400 58.805 21.660 59.065 ;
        RECT 21.400 58.145 21.660 58.405 ;
        RECT 21.400 57.485 21.660 57.745 ;
        RECT 21.400 56.825 21.660 57.085 ;
        RECT 21.400 56.165 21.660 56.425 ;
        RECT 21.400 55.505 21.660 55.765 ;
        RECT 21.400 54.845 21.660 55.105 ;
        RECT 21.400 54.185 21.660 54.445 ;
        RECT 21.400 53.525 21.660 53.785 ;
        RECT 21.400 52.865 21.660 53.125 ;
        RECT 21.400 52.205 21.660 52.465 ;
        RECT 21.400 51.545 21.660 51.805 ;
        RECT 21.400 50.885 21.660 51.145 ;
        RECT 21.400 50.225 21.660 50.485 ;
        RECT 25.885 42.465 26.145 42.725 ;
        RECT 26.545 42.465 26.805 42.725 ;
        RECT 27.205 42.465 27.465 42.725 ;
        RECT 25.885 41.805 26.145 42.065 ;
        RECT 26.545 41.805 26.805 42.065 ;
        RECT 27.205 41.805 27.465 42.065 ;
        RECT 25.885 41.145 26.145 41.405 ;
        RECT 26.545 41.145 26.805 41.405 ;
        RECT 27.205 41.145 27.465 41.405 ;
        RECT 25.885 27.665 26.145 27.925 ;
        RECT 26.545 27.665 26.805 27.925 ;
        RECT 27.205 27.665 27.465 27.925 ;
        RECT 25.885 27.005 26.145 27.265 ;
        RECT 26.545 27.005 26.805 27.265 ;
        RECT 27.205 27.005 27.465 27.265 ;
        RECT 25.885 26.345 26.145 26.605 ;
        RECT 26.545 26.345 26.805 26.605 ;
        RECT 27.205 26.345 27.465 26.605 ;
        RECT 31.690 58.805 31.950 59.065 ;
        RECT 31.690 58.145 31.950 58.405 ;
        RECT 31.690 57.485 31.950 57.745 ;
        RECT 31.690 56.825 31.950 57.085 ;
        RECT 31.690 56.165 31.950 56.425 ;
        RECT 31.690 55.505 31.950 55.765 ;
        RECT 31.690 54.845 31.950 55.105 ;
        RECT 31.690 54.185 31.950 54.445 ;
        RECT 31.690 53.525 31.950 53.785 ;
        RECT 31.690 52.865 31.950 53.125 ;
        RECT 31.690 52.205 31.950 52.465 ;
        RECT 31.690 51.545 31.950 51.805 ;
        RECT 31.690 50.885 31.950 51.145 ;
        RECT 31.690 50.225 31.950 50.485 ;
        RECT 44.760 59.990 45.020 60.250 ;
        RECT 62.605 59.990 62.865 60.250 ;
        RECT 36.185 39.765 36.445 40.025 ;
        RECT 36.845 39.765 37.105 40.025 ;
        RECT 37.505 39.765 37.765 40.025 ;
        RECT 36.185 39.105 36.445 39.365 ;
        RECT 36.845 39.105 37.105 39.365 ;
        RECT 37.505 39.105 37.765 39.365 ;
        RECT 36.185 38.445 36.445 38.705 ;
        RECT 36.845 38.445 37.105 38.705 ;
        RECT 37.505 38.445 37.765 38.705 ;
        RECT 36.185 30.365 36.445 30.625 ;
        RECT 36.845 30.365 37.105 30.625 ;
        RECT 37.505 30.365 37.765 30.625 ;
        RECT 36.185 29.705 36.445 29.965 ;
        RECT 36.845 29.705 37.105 29.965 ;
        RECT 37.505 29.705 37.765 29.965 ;
        RECT 36.185 29.045 36.445 29.305 ;
        RECT 36.845 29.045 37.105 29.305 ;
        RECT 37.505 29.045 37.765 29.305 ;
        RECT 12.480 8.805 12.740 9.065 ;
        RECT 30.325 8.805 30.585 9.065 ;
        RECT 41.975 58.805 42.235 59.065 ;
        RECT 41.975 58.145 42.235 58.405 ;
        RECT 41.975 57.485 42.235 57.745 ;
        RECT 41.975 56.825 42.235 57.085 ;
        RECT 41.975 56.165 42.235 56.425 ;
        RECT 41.975 55.505 42.235 55.765 ;
        RECT 41.975 54.845 42.235 55.105 ;
        RECT 41.975 54.185 42.235 54.445 ;
        RECT 41.975 53.525 42.235 53.785 ;
        RECT 41.975 52.865 42.235 53.125 ;
        RECT 41.975 52.205 42.235 52.465 ;
        RECT 41.975 51.545 42.235 51.805 ;
        RECT 41.975 50.885 42.235 51.145 ;
        RECT 41.975 50.225 42.235 50.485 ;
        RECT 43.395 58.805 43.655 59.065 ;
        RECT 43.395 58.145 43.655 58.405 ;
        RECT 43.395 57.485 43.655 57.745 ;
        RECT 43.395 56.825 43.655 57.085 ;
        RECT 43.395 56.165 43.655 56.425 ;
        RECT 43.395 55.505 43.655 55.765 ;
        RECT 43.395 54.845 43.655 55.105 ;
        RECT 43.395 54.185 43.655 54.445 ;
        RECT 43.395 53.525 43.655 53.785 ;
        RECT 43.395 52.865 43.655 53.125 ;
        RECT 43.395 52.205 43.655 52.465 ;
        RECT 43.395 51.545 43.655 51.805 ;
        RECT 43.395 50.885 43.655 51.145 ;
        RECT 43.395 50.225 43.655 50.485 ;
        RECT 47.880 47.865 48.140 48.125 ;
        RECT 48.540 47.865 48.800 48.125 ;
        RECT 49.200 47.865 49.460 48.125 ;
        RECT 47.880 47.205 48.140 47.465 ;
        RECT 48.540 47.205 48.800 47.465 ;
        RECT 49.200 47.205 49.460 47.465 ;
        RECT 47.880 46.545 48.140 46.805 ;
        RECT 48.540 46.545 48.800 46.805 ;
        RECT 49.200 46.545 49.460 46.805 ;
        RECT 47.880 22.265 48.140 22.525 ;
        RECT 48.540 22.265 48.800 22.525 ;
        RECT 49.200 22.265 49.460 22.525 ;
        RECT 47.880 21.605 48.140 21.865 ;
        RECT 48.540 21.605 48.800 21.865 ;
        RECT 49.200 21.605 49.460 21.865 ;
        RECT 47.880 20.945 48.140 21.205 ;
        RECT 48.540 20.945 48.800 21.205 ;
        RECT 49.200 20.945 49.460 21.205 ;
        RECT 53.685 58.805 53.945 59.065 ;
        RECT 53.685 58.145 53.945 58.405 ;
        RECT 53.685 57.485 53.945 57.745 ;
        RECT 53.685 56.825 53.945 57.085 ;
        RECT 53.685 56.165 53.945 56.425 ;
        RECT 53.685 55.505 53.945 55.765 ;
        RECT 53.685 54.845 53.945 55.105 ;
        RECT 53.685 54.185 53.945 54.445 ;
        RECT 53.685 53.525 53.945 53.785 ;
        RECT 53.685 52.865 53.945 53.125 ;
        RECT 53.685 52.205 53.945 52.465 ;
        RECT 53.685 51.545 53.945 51.805 ;
        RECT 53.685 50.885 53.945 51.145 ;
        RECT 53.685 50.225 53.945 50.485 ;
        RECT 65.335 59.990 65.595 60.250 ;
        RECT 83.180 59.990 83.440 60.250 ;
        RECT 58.180 45.165 58.440 45.425 ;
        RECT 58.840 45.165 59.100 45.425 ;
        RECT 59.500 45.165 59.760 45.425 ;
        RECT 58.180 44.505 58.440 44.765 ;
        RECT 58.840 44.505 59.100 44.765 ;
        RECT 59.500 44.505 59.760 44.765 ;
        RECT 58.180 43.845 58.440 44.105 ;
        RECT 58.840 43.845 59.100 44.105 ;
        RECT 59.500 43.845 59.760 44.105 ;
        RECT 58.180 24.965 58.440 25.225 ;
        RECT 58.840 24.965 59.100 25.225 ;
        RECT 59.500 24.965 59.760 25.225 ;
        RECT 58.180 24.305 58.440 24.565 ;
        RECT 58.840 24.305 59.100 24.565 ;
        RECT 59.500 24.305 59.760 24.565 ;
        RECT 58.180 23.645 58.440 23.905 ;
        RECT 58.840 23.645 59.100 23.905 ;
        RECT 59.500 23.645 59.760 23.905 ;
        RECT 33.055 8.805 33.315 9.065 ;
        RECT 52.320 8.805 52.580 9.065 ;
        RECT 63.970 58.805 64.230 59.065 ;
        RECT 63.970 58.145 64.230 58.405 ;
        RECT 63.970 57.485 64.230 57.745 ;
        RECT 63.970 56.825 64.230 57.085 ;
        RECT 63.970 56.165 64.230 56.425 ;
        RECT 63.970 55.505 64.230 55.765 ;
        RECT 63.970 54.845 64.230 55.105 ;
        RECT 63.970 54.185 64.230 54.445 ;
        RECT 63.970 53.525 64.230 53.785 ;
        RECT 63.970 52.865 64.230 53.125 ;
        RECT 63.970 52.205 64.230 52.465 ;
        RECT 63.970 51.545 64.230 51.805 ;
        RECT 63.970 50.885 64.230 51.145 ;
        RECT 63.970 50.225 64.230 50.485 ;
        RECT 68.455 42.465 68.715 42.725 ;
        RECT 69.115 42.465 69.375 42.725 ;
        RECT 69.775 42.465 70.035 42.725 ;
        RECT 68.455 41.805 68.715 42.065 ;
        RECT 69.115 41.805 69.375 42.065 ;
        RECT 69.775 41.805 70.035 42.065 ;
        RECT 68.455 41.145 68.715 41.405 ;
        RECT 69.115 41.145 69.375 41.405 ;
        RECT 69.775 41.145 70.035 41.405 ;
        RECT 68.455 27.665 68.715 27.925 ;
        RECT 69.115 27.665 69.375 27.925 ;
        RECT 69.775 27.665 70.035 27.925 ;
        RECT 68.455 27.005 68.715 27.265 ;
        RECT 69.115 27.005 69.375 27.265 ;
        RECT 69.775 27.005 70.035 27.265 ;
        RECT 68.455 26.345 68.715 26.605 ;
        RECT 69.115 26.345 69.375 26.605 ;
        RECT 69.775 26.345 70.035 26.605 ;
        RECT 74.260 58.805 74.520 59.065 ;
        RECT 74.260 58.145 74.520 58.405 ;
        RECT 74.260 57.485 74.520 57.745 ;
        RECT 74.260 56.825 74.520 57.085 ;
        RECT 74.260 56.165 74.520 56.425 ;
        RECT 74.260 55.505 74.520 55.765 ;
        RECT 74.260 54.845 74.520 55.105 ;
        RECT 74.260 54.185 74.520 54.445 ;
        RECT 74.260 53.525 74.520 53.785 ;
        RECT 74.260 52.865 74.520 53.125 ;
        RECT 74.260 52.205 74.520 52.465 ;
        RECT 74.260 51.545 74.520 51.805 ;
        RECT 74.260 50.885 74.520 51.145 ;
        RECT 74.260 50.225 74.520 50.485 ;
        RECT 87.330 59.990 87.590 60.250 ;
        RECT 105.175 59.990 105.435 60.250 ;
        RECT 78.755 39.765 79.015 40.025 ;
        RECT 79.415 39.765 79.675 40.025 ;
        RECT 80.075 39.765 80.335 40.025 ;
        RECT 78.755 39.105 79.015 39.365 ;
        RECT 79.415 39.105 79.675 39.365 ;
        RECT 80.075 39.105 80.335 39.365 ;
        RECT 78.755 38.445 79.015 38.705 ;
        RECT 79.415 38.445 79.675 38.705 ;
        RECT 80.075 38.445 80.335 38.705 ;
        RECT 78.755 30.365 79.015 30.625 ;
        RECT 79.415 30.365 79.675 30.625 ;
        RECT 80.075 30.365 80.335 30.625 ;
        RECT 78.755 29.705 79.015 29.965 ;
        RECT 79.415 29.705 79.675 29.965 ;
        RECT 80.075 29.705 80.335 29.965 ;
        RECT 78.755 29.045 79.015 29.305 ;
        RECT 79.415 29.045 79.675 29.305 ;
        RECT 80.075 29.045 80.335 29.305 ;
        RECT 55.050 8.805 55.310 9.065 ;
        RECT 72.895 8.805 73.155 9.065 ;
        RECT 84.545 58.805 84.805 59.065 ;
        RECT 84.545 58.145 84.805 58.405 ;
        RECT 84.545 57.485 84.805 57.745 ;
        RECT 84.545 56.825 84.805 57.085 ;
        RECT 84.545 56.165 84.805 56.425 ;
        RECT 84.545 55.505 84.805 55.765 ;
        RECT 84.545 54.845 84.805 55.105 ;
        RECT 84.545 54.185 84.805 54.445 ;
        RECT 84.545 53.525 84.805 53.785 ;
        RECT 84.545 52.865 84.805 53.125 ;
        RECT 84.545 52.205 84.805 52.465 ;
        RECT 84.545 51.545 84.805 51.805 ;
        RECT 84.545 50.885 84.805 51.145 ;
        RECT 84.545 50.225 84.805 50.485 ;
        RECT 85.965 58.805 86.225 59.065 ;
        RECT 85.965 58.145 86.225 58.405 ;
        RECT 85.965 57.485 86.225 57.745 ;
        RECT 85.965 56.825 86.225 57.085 ;
        RECT 85.965 56.165 86.225 56.425 ;
        RECT 85.965 55.505 86.225 55.765 ;
        RECT 85.965 54.845 86.225 55.105 ;
        RECT 85.965 54.185 86.225 54.445 ;
        RECT 85.965 53.525 86.225 53.785 ;
        RECT 85.965 52.865 86.225 53.125 ;
        RECT 85.965 52.205 86.225 52.465 ;
        RECT 85.965 51.545 86.225 51.805 ;
        RECT 85.965 50.885 86.225 51.145 ;
        RECT 85.965 50.225 86.225 50.485 ;
        RECT 90.450 47.865 90.710 48.125 ;
        RECT 91.110 47.865 91.370 48.125 ;
        RECT 91.770 47.865 92.030 48.125 ;
        RECT 90.450 47.205 90.710 47.465 ;
        RECT 91.110 47.205 91.370 47.465 ;
        RECT 91.770 47.205 92.030 47.465 ;
        RECT 90.450 46.545 90.710 46.805 ;
        RECT 91.110 46.545 91.370 46.805 ;
        RECT 91.770 46.545 92.030 46.805 ;
        RECT 90.450 22.265 90.710 22.525 ;
        RECT 91.110 22.265 91.370 22.525 ;
        RECT 91.770 22.265 92.030 22.525 ;
        RECT 90.450 21.605 90.710 21.865 ;
        RECT 91.110 21.605 91.370 21.865 ;
        RECT 91.770 21.605 92.030 21.865 ;
        RECT 90.450 20.945 90.710 21.205 ;
        RECT 91.110 20.945 91.370 21.205 ;
        RECT 91.770 20.945 92.030 21.205 ;
        RECT 96.255 58.805 96.515 59.065 ;
        RECT 96.255 58.145 96.515 58.405 ;
        RECT 96.255 57.485 96.515 57.745 ;
        RECT 96.255 56.825 96.515 57.085 ;
        RECT 96.255 56.165 96.515 56.425 ;
        RECT 96.255 55.505 96.515 55.765 ;
        RECT 96.255 54.845 96.515 55.105 ;
        RECT 96.255 54.185 96.515 54.445 ;
        RECT 96.255 53.525 96.515 53.785 ;
        RECT 96.255 52.865 96.515 53.125 ;
        RECT 96.255 52.205 96.515 52.465 ;
        RECT 96.255 51.545 96.515 51.805 ;
        RECT 96.255 50.885 96.515 51.145 ;
        RECT 96.255 50.225 96.515 50.485 ;
        RECT 107.905 59.990 108.165 60.250 ;
        RECT 125.750 59.990 126.010 60.250 ;
        RECT 100.750 45.165 101.010 45.425 ;
        RECT 101.410 45.165 101.670 45.425 ;
        RECT 102.070 45.165 102.330 45.425 ;
        RECT 100.750 44.505 101.010 44.765 ;
        RECT 101.410 44.505 101.670 44.765 ;
        RECT 102.070 44.505 102.330 44.765 ;
        RECT 100.750 43.845 101.010 44.105 ;
        RECT 101.410 43.845 101.670 44.105 ;
        RECT 102.070 43.845 102.330 44.105 ;
        RECT 100.750 24.965 101.010 25.225 ;
        RECT 101.410 24.965 101.670 25.225 ;
        RECT 102.070 24.965 102.330 25.225 ;
        RECT 100.750 24.305 101.010 24.565 ;
        RECT 101.410 24.305 101.670 24.565 ;
        RECT 102.070 24.305 102.330 24.565 ;
        RECT 100.750 23.645 101.010 23.905 ;
        RECT 101.410 23.645 101.670 23.905 ;
        RECT 102.070 23.645 102.330 23.905 ;
        RECT 75.625 8.805 75.885 9.065 ;
        RECT 94.890 8.805 95.150 9.065 ;
        RECT 106.540 58.805 106.800 59.065 ;
        RECT 106.540 58.145 106.800 58.405 ;
        RECT 106.540 57.485 106.800 57.745 ;
        RECT 106.540 56.825 106.800 57.085 ;
        RECT 106.540 56.165 106.800 56.425 ;
        RECT 106.540 55.505 106.800 55.765 ;
        RECT 106.540 54.845 106.800 55.105 ;
        RECT 106.540 54.185 106.800 54.445 ;
        RECT 106.540 53.525 106.800 53.785 ;
        RECT 106.540 52.865 106.800 53.125 ;
        RECT 106.540 52.205 106.800 52.465 ;
        RECT 106.540 51.545 106.800 51.805 ;
        RECT 106.540 50.885 106.800 51.145 ;
        RECT 106.540 50.225 106.800 50.485 ;
        RECT 111.025 42.465 111.285 42.725 ;
        RECT 111.685 42.465 111.945 42.725 ;
        RECT 112.345 42.465 112.605 42.725 ;
        RECT 111.025 41.805 111.285 42.065 ;
        RECT 111.685 41.805 111.945 42.065 ;
        RECT 112.345 41.805 112.605 42.065 ;
        RECT 111.025 41.145 111.285 41.405 ;
        RECT 111.685 41.145 111.945 41.405 ;
        RECT 112.345 41.145 112.605 41.405 ;
        RECT 111.025 27.665 111.285 27.925 ;
        RECT 111.685 27.665 111.945 27.925 ;
        RECT 112.345 27.665 112.605 27.925 ;
        RECT 111.025 27.005 111.285 27.265 ;
        RECT 111.685 27.005 111.945 27.265 ;
        RECT 112.345 27.005 112.605 27.265 ;
        RECT 111.025 26.345 111.285 26.605 ;
        RECT 111.685 26.345 111.945 26.605 ;
        RECT 112.345 26.345 112.605 26.605 ;
        RECT 116.830 58.805 117.090 59.065 ;
        RECT 116.830 58.145 117.090 58.405 ;
        RECT 116.830 57.485 117.090 57.745 ;
        RECT 116.830 56.825 117.090 57.085 ;
        RECT 116.830 56.165 117.090 56.425 ;
        RECT 116.830 55.505 117.090 55.765 ;
        RECT 116.830 54.845 117.090 55.105 ;
        RECT 116.830 54.185 117.090 54.445 ;
        RECT 116.830 53.525 117.090 53.785 ;
        RECT 116.830 52.865 117.090 53.125 ;
        RECT 116.830 52.205 117.090 52.465 ;
        RECT 116.830 51.545 117.090 51.805 ;
        RECT 116.830 50.885 117.090 51.145 ;
        RECT 116.830 50.225 117.090 50.485 ;
        RECT 129.900 59.990 130.160 60.250 ;
        RECT 147.745 59.990 148.005 60.250 ;
        RECT 121.325 39.765 121.585 40.025 ;
        RECT 121.985 39.765 122.245 40.025 ;
        RECT 122.645 39.765 122.905 40.025 ;
        RECT 121.325 39.105 121.585 39.365 ;
        RECT 121.985 39.105 122.245 39.365 ;
        RECT 122.645 39.105 122.905 39.365 ;
        RECT 121.325 38.445 121.585 38.705 ;
        RECT 121.985 38.445 122.245 38.705 ;
        RECT 122.645 38.445 122.905 38.705 ;
        RECT 121.325 30.365 121.585 30.625 ;
        RECT 121.985 30.365 122.245 30.625 ;
        RECT 122.645 30.365 122.905 30.625 ;
        RECT 121.325 29.705 121.585 29.965 ;
        RECT 121.985 29.705 122.245 29.965 ;
        RECT 122.645 29.705 122.905 29.965 ;
        RECT 121.325 29.045 121.585 29.305 ;
        RECT 121.985 29.045 122.245 29.305 ;
        RECT 122.645 29.045 122.905 29.305 ;
        RECT 97.620 8.805 97.880 9.065 ;
        RECT 115.465 8.805 115.725 9.065 ;
        RECT 127.115 58.805 127.375 59.065 ;
        RECT 127.115 58.145 127.375 58.405 ;
        RECT 127.115 57.485 127.375 57.745 ;
        RECT 127.115 56.825 127.375 57.085 ;
        RECT 127.115 56.165 127.375 56.425 ;
        RECT 127.115 55.505 127.375 55.765 ;
        RECT 127.115 54.845 127.375 55.105 ;
        RECT 127.115 54.185 127.375 54.445 ;
        RECT 127.115 53.525 127.375 53.785 ;
        RECT 127.115 52.865 127.375 53.125 ;
        RECT 127.115 52.205 127.375 52.465 ;
        RECT 127.115 51.545 127.375 51.805 ;
        RECT 127.115 50.885 127.375 51.145 ;
        RECT 127.115 50.225 127.375 50.485 ;
        RECT 128.535 58.805 128.795 59.065 ;
        RECT 128.535 58.145 128.795 58.405 ;
        RECT 128.535 57.485 128.795 57.745 ;
        RECT 128.535 56.825 128.795 57.085 ;
        RECT 128.535 56.165 128.795 56.425 ;
        RECT 128.535 55.505 128.795 55.765 ;
        RECT 128.535 54.845 128.795 55.105 ;
        RECT 128.535 54.185 128.795 54.445 ;
        RECT 128.535 53.525 128.795 53.785 ;
        RECT 128.535 52.865 128.795 53.125 ;
        RECT 128.535 52.205 128.795 52.465 ;
        RECT 128.535 51.545 128.795 51.805 ;
        RECT 128.535 50.885 128.795 51.145 ;
        RECT 128.535 50.225 128.795 50.485 ;
        RECT 133.020 47.865 133.280 48.125 ;
        RECT 133.680 47.865 133.940 48.125 ;
        RECT 134.340 47.865 134.600 48.125 ;
        RECT 133.020 47.205 133.280 47.465 ;
        RECT 133.680 47.205 133.940 47.465 ;
        RECT 134.340 47.205 134.600 47.465 ;
        RECT 133.020 46.545 133.280 46.805 ;
        RECT 133.680 46.545 133.940 46.805 ;
        RECT 134.340 46.545 134.600 46.805 ;
        RECT 133.020 22.265 133.280 22.525 ;
        RECT 133.680 22.265 133.940 22.525 ;
        RECT 134.340 22.265 134.600 22.525 ;
        RECT 133.020 21.605 133.280 21.865 ;
        RECT 133.680 21.605 133.940 21.865 ;
        RECT 134.340 21.605 134.600 21.865 ;
        RECT 133.020 20.945 133.280 21.205 ;
        RECT 133.680 20.945 133.940 21.205 ;
        RECT 134.340 20.945 134.600 21.205 ;
        RECT 138.825 58.805 139.085 59.065 ;
        RECT 138.825 58.145 139.085 58.405 ;
        RECT 138.825 57.485 139.085 57.745 ;
        RECT 138.825 56.825 139.085 57.085 ;
        RECT 138.825 56.165 139.085 56.425 ;
        RECT 138.825 55.505 139.085 55.765 ;
        RECT 138.825 54.845 139.085 55.105 ;
        RECT 138.825 54.185 139.085 54.445 ;
        RECT 138.825 53.525 139.085 53.785 ;
        RECT 138.825 52.865 139.085 53.125 ;
        RECT 138.825 52.205 139.085 52.465 ;
        RECT 138.825 51.545 139.085 51.805 ;
        RECT 138.825 50.885 139.085 51.145 ;
        RECT 138.825 50.225 139.085 50.485 ;
        RECT 150.475 59.990 150.735 60.250 ;
        RECT 168.320 59.990 168.580 60.250 ;
        RECT 143.320 45.165 143.580 45.425 ;
        RECT 143.980 45.165 144.240 45.425 ;
        RECT 144.640 45.165 144.900 45.425 ;
        RECT 143.320 44.505 143.580 44.765 ;
        RECT 143.980 44.505 144.240 44.765 ;
        RECT 144.640 44.505 144.900 44.765 ;
        RECT 143.320 43.845 143.580 44.105 ;
        RECT 143.980 43.845 144.240 44.105 ;
        RECT 144.640 43.845 144.900 44.105 ;
        RECT 143.320 24.965 143.580 25.225 ;
        RECT 143.980 24.965 144.240 25.225 ;
        RECT 144.640 24.965 144.900 25.225 ;
        RECT 143.320 24.305 143.580 24.565 ;
        RECT 143.980 24.305 144.240 24.565 ;
        RECT 144.640 24.305 144.900 24.565 ;
        RECT 143.320 23.645 143.580 23.905 ;
        RECT 143.980 23.645 144.240 23.905 ;
        RECT 144.640 23.645 144.900 23.905 ;
        RECT 118.195 8.805 118.455 9.065 ;
        RECT 137.460 8.805 137.720 9.065 ;
        RECT 149.110 58.805 149.370 59.065 ;
        RECT 149.110 58.145 149.370 58.405 ;
        RECT 149.110 57.485 149.370 57.745 ;
        RECT 149.110 56.825 149.370 57.085 ;
        RECT 149.110 56.165 149.370 56.425 ;
        RECT 149.110 55.505 149.370 55.765 ;
        RECT 149.110 54.845 149.370 55.105 ;
        RECT 149.110 54.185 149.370 54.445 ;
        RECT 149.110 53.525 149.370 53.785 ;
        RECT 149.110 52.865 149.370 53.125 ;
        RECT 149.110 52.205 149.370 52.465 ;
        RECT 149.110 51.545 149.370 51.805 ;
        RECT 149.110 50.885 149.370 51.145 ;
        RECT 149.110 50.225 149.370 50.485 ;
        RECT 153.595 42.465 153.855 42.725 ;
        RECT 154.255 42.465 154.515 42.725 ;
        RECT 154.915 42.465 155.175 42.725 ;
        RECT 153.595 41.805 153.855 42.065 ;
        RECT 154.255 41.805 154.515 42.065 ;
        RECT 154.915 41.805 155.175 42.065 ;
        RECT 153.595 41.145 153.855 41.405 ;
        RECT 154.255 41.145 154.515 41.405 ;
        RECT 154.915 41.145 155.175 41.405 ;
        RECT 153.595 27.665 153.855 27.925 ;
        RECT 154.255 27.665 154.515 27.925 ;
        RECT 154.915 27.665 155.175 27.925 ;
        RECT 153.595 27.005 153.855 27.265 ;
        RECT 154.255 27.005 154.515 27.265 ;
        RECT 154.915 27.005 155.175 27.265 ;
        RECT 153.595 26.345 153.855 26.605 ;
        RECT 154.255 26.345 154.515 26.605 ;
        RECT 154.915 26.345 155.175 26.605 ;
        RECT 159.400 58.805 159.660 59.065 ;
        RECT 159.400 58.145 159.660 58.405 ;
        RECT 159.400 57.485 159.660 57.745 ;
        RECT 159.400 56.825 159.660 57.085 ;
        RECT 159.400 56.165 159.660 56.425 ;
        RECT 159.400 55.505 159.660 55.765 ;
        RECT 159.400 54.845 159.660 55.105 ;
        RECT 159.400 54.185 159.660 54.445 ;
        RECT 159.400 53.525 159.660 53.785 ;
        RECT 159.400 52.865 159.660 53.125 ;
        RECT 159.400 52.205 159.660 52.465 ;
        RECT 159.400 51.545 159.660 51.805 ;
        RECT 159.400 50.885 159.660 51.145 ;
        RECT 159.400 50.225 159.660 50.485 ;
        RECT 172.470 59.990 172.730 60.250 ;
        RECT 190.315 59.990 190.575 60.250 ;
        RECT 163.895 39.765 164.155 40.025 ;
        RECT 164.555 39.765 164.815 40.025 ;
        RECT 165.215 39.765 165.475 40.025 ;
        RECT 163.895 39.105 164.155 39.365 ;
        RECT 164.555 39.105 164.815 39.365 ;
        RECT 165.215 39.105 165.475 39.365 ;
        RECT 163.895 38.445 164.155 38.705 ;
        RECT 164.555 38.445 164.815 38.705 ;
        RECT 165.215 38.445 165.475 38.705 ;
        RECT 163.895 30.365 164.155 30.625 ;
        RECT 164.555 30.365 164.815 30.625 ;
        RECT 165.215 30.365 165.475 30.625 ;
        RECT 163.895 29.705 164.155 29.965 ;
        RECT 164.555 29.705 164.815 29.965 ;
        RECT 165.215 29.705 165.475 29.965 ;
        RECT 163.895 29.045 164.155 29.305 ;
        RECT 164.555 29.045 164.815 29.305 ;
        RECT 165.215 29.045 165.475 29.305 ;
        RECT 140.190 8.805 140.450 9.065 ;
        RECT 158.035 8.805 158.295 9.065 ;
        RECT 169.685 58.805 169.945 59.065 ;
        RECT 169.685 58.145 169.945 58.405 ;
        RECT 169.685 57.485 169.945 57.745 ;
        RECT 169.685 56.825 169.945 57.085 ;
        RECT 169.685 56.165 169.945 56.425 ;
        RECT 169.685 55.505 169.945 55.765 ;
        RECT 169.685 54.845 169.945 55.105 ;
        RECT 169.685 54.185 169.945 54.445 ;
        RECT 169.685 53.525 169.945 53.785 ;
        RECT 169.685 52.865 169.945 53.125 ;
        RECT 169.685 52.205 169.945 52.465 ;
        RECT 169.685 51.545 169.945 51.805 ;
        RECT 169.685 50.885 169.945 51.145 ;
        RECT 169.685 50.225 169.945 50.485 ;
        RECT 171.105 58.805 171.365 59.065 ;
        RECT 171.105 58.145 171.365 58.405 ;
        RECT 171.105 57.485 171.365 57.745 ;
        RECT 171.105 56.825 171.365 57.085 ;
        RECT 171.105 56.165 171.365 56.425 ;
        RECT 171.105 55.505 171.365 55.765 ;
        RECT 171.105 54.845 171.365 55.105 ;
        RECT 171.105 54.185 171.365 54.445 ;
        RECT 171.105 53.525 171.365 53.785 ;
        RECT 171.105 52.865 171.365 53.125 ;
        RECT 171.105 52.205 171.365 52.465 ;
        RECT 171.105 51.545 171.365 51.805 ;
        RECT 171.105 50.885 171.365 51.145 ;
        RECT 171.105 50.225 171.365 50.485 ;
        RECT 175.590 47.865 175.850 48.125 ;
        RECT 176.250 47.865 176.510 48.125 ;
        RECT 176.910 47.865 177.170 48.125 ;
        RECT 175.590 47.205 175.850 47.465 ;
        RECT 176.250 47.205 176.510 47.465 ;
        RECT 176.910 47.205 177.170 47.465 ;
        RECT 175.590 46.545 175.850 46.805 ;
        RECT 176.250 46.545 176.510 46.805 ;
        RECT 176.910 46.545 177.170 46.805 ;
        RECT 175.590 22.265 175.850 22.525 ;
        RECT 176.250 22.265 176.510 22.525 ;
        RECT 176.910 22.265 177.170 22.525 ;
        RECT 175.590 21.605 175.850 21.865 ;
        RECT 176.250 21.605 176.510 21.865 ;
        RECT 176.910 21.605 177.170 21.865 ;
        RECT 175.590 20.945 175.850 21.205 ;
        RECT 176.250 20.945 176.510 21.205 ;
        RECT 176.910 20.945 177.170 21.205 ;
        RECT 181.395 58.805 181.655 59.065 ;
        RECT 181.395 58.145 181.655 58.405 ;
        RECT 181.395 57.485 181.655 57.745 ;
        RECT 181.395 56.825 181.655 57.085 ;
        RECT 181.395 56.165 181.655 56.425 ;
        RECT 181.395 55.505 181.655 55.765 ;
        RECT 181.395 54.845 181.655 55.105 ;
        RECT 181.395 54.185 181.655 54.445 ;
        RECT 181.395 53.525 181.655 53.785 ;
        RECT 181.395 52.865 181.655 53.125 ;
        RECT 181.395 52.205 181.655 52.465 ;
        RECT 181.395 51.545 181.655 51.805 ;
        RECT 181.395 50.885 181.655 51.145 ;
        RECT 181.395 50.225 181.655 50.485 ;
        RECT 193.045 59.990 193.305 60.250 ;
        RECT 210.890 59.990 211.150 60.250 ;
        RECT 185.890 45.165 186.150 45.425 ;
        RECT 186.550 45.165 186.810 45.425 ;
        RECT 187.210 45.165 187.470 45.425 ;
        RECT 185.890 44.505 186.150 44.765 ;
        RECT 186.550 44.505 186.810 44.765 ;
        RECT 187.210 44.505 187.470 44.765 ;
        RECT 185.890 43.845 186.150 44.105 ;
        RECT 186.550 43.845 186.810 44.105 ;
        RECT 187.210 43.845 187.470 44.105 ;
        RECT 185.890 24.965 186.150 25.225 ;
        RECT 186.550 24.965 186.810 25.225 ;
        RECT 187.210 24.965 187.470 25.225 ;
        RECT 185.890 24.305 186.150 24.565 ;
        RECT 186.550 24.305 186.810 24.565 ;
        RECT 187.210 24.305 187.470 24.565 ;
        RECT 185.890 23.645 186.150 23.905 ;
        RECT 186.550 23.645 186.810 23.905 ;
        RECT 187.210 23.645 187.470 23.905 ;
        RECT 160.765 8.805 161.025 9.065 ;
        RECT 180.030 8.805 180.290 9.065 ;
        RECT 191.680 58.805 191.940 59.065 ;
        RECT 191.680 58.145 191.940 58.405 ;
        RECT 191.680 57.485 191.940 57.745 ;
        RECT 191.680 56.825 191.940 57.085 ;
        RECT 191.680 56.165 191.940 56.425 ;
        RECT 191.680 55.505 191.940 55.765 ;
        RECT 191.680 54.845 191.940 55.105 ;
        RECT 191.680 54.185 191.940 54.445 ;
        RECT 191.680 53.525 191.940 53.785 ;
        RECT 191.680 52.865 191.940 53.125 ;
        RECT 191.680 52.205 191.940 52.465 ;
        RECT 191.680 51.545 191.940 51.805 ;
        RECT 191.680 50.885 191.940 51.145 ;
        RECT 191.680 50.225 191.940 50.485 ;
        RECT 196.165 42.465 196.425 42.725 ;
        RECT 196.825 42.465 197.085 42.725 ;
        RECT 197.485 42.465 197.745 42.725 ;
        RECT 196.165 41.805 196.425 42.065 ;
        RECT 196.825 41.805 197.085 42.065 ;
        RECT 197.485 41.805 197.745 42.065 ;
        RECT 196.165 41.145 196.425 41.405 ;
        RECT 196.825 41.145 197.085 41.405 ;
        RECT 197.485 41.145 197.745 41.405 ;
        RECT 196.165 27.665 196.425 27.925 ;
        RECT 196.825 27.665 197.085 27.925 ;
        RECT 197.485 27.665 197.745 27.925 ;
        RECT 196.165 27.005 196.425 27.265 ;
        RECT 196.825 27.005 197.085 27.265 ;
        RECT 197.485 27.005 197.745 27.265 ;
        RECT 196.165 26.345 196.425 26.605 ;
        RECT 196.825 26.345 197.085 26.605 ;
        RECT 197.485 26.345 197.745 26.605 ;
        RECT 201.970 58.805 202.230 59.065 ;
        RECT 201.970 58.145 202.230 58.405 ;
        RECT 201.970 57.485 202.230 57.745 ;
        RECT 201.970 56.825 202.230 57.085 ;
        RECT 201.970 56.165 202.230 56.425 ;
        RECT 201.970 55.505 202.230 55.765 ;
        RECT 201.970 54.845 202.230 55.105 ;
        RECT 201.970 54.185 202.230 54.445 ;
        RECT 201.970 53.525 202.230 53.785 ;
        RECT 201.970 52.865 202.230 53.125 ;
        RECT 201.970 52.205 202.230 52.465 ;
        RECT 201.970 51.545 202.230 51.805 ;
        RECT 201.970 50.885 202.230 51.145 ;
        RECT 201.970 50.225 202.230 50.485 ;
        RECT 215.040 59.990 215.300 60.250 ;
        RECT 232.885 59.990 233.145 60.250 ;
        RECT 206.465 39.765 206.725 40.025 ;
        RECT 207.125 39.765 207.385 40.025 ;
        RECT 207.785 39.765 208.045 40.025 ;
        RECT 206.465 39.105 206.725 39.365 ;
        RECT 207.125 39.105 207.385 39.365 ;
        RECT 207.785 39.105 208.045 39.365 ;
        RECT 206.465 38.445 206.725 38.705 ;
        RECT 207.125 38.445 207.385 38.705 ;
        RECT 207.785 38.445 208.045 38.705 ;
        RECT 206.465 30.365 206.725 30.625 ;
        RECT 207.125 30.365 207.385 30.625 ;
        RECT 207.785 30.365 208.045 30.625 ;
        RECT 206.465 29.705 206.725 29.965 ;
        RECT 207.125 29.705 207.385 29.965 ;
        RECT 207.785 29.705 208.045 29.965 ;
        RECT 206.465 29.045 206.725 29.305 ;
        RECT 207.125 29.045 207.385 29.305 ;
        RECT 207.785 29.045 208.045 29.305 ;
        RECT 182.760 8.805 183.020 9.065 ;
        RECT 200.605 8.805 200.865 9.065 ;
        RECT 212.255 58.805 212.515 59.065 ;
        RECT 212.255 58.145 212.515 58.405 ;
        RECT 212.255 57.485 212.515 57.745 ;
        RECT 212.255 56.825 212.515 57.085 ;
        RECT 212.255 56.165 212.515 56.425 ;
        RECT 212.255 55.505 212.515 55.765 ;
        RECT 212.255 54.845 212.515 55.105 ;
        RECT 212.255 54.185 212.515 54.445 ;
        RECT 212.255 53.525 212.515 53.785 ;
        RECT 212.255 52.865 212.515 53.125 ;
        RECT 212.255 52.205 212.515 52.465 ;
        RECT 212.255 51.545 212.515 51.805 ;
        RECT 212.255 50.885 212.515 51.145 ;
        RECT 212.255 50.225 212.515 50.485 ;
        RECT 213.675 58.805 213.935 59.065 ;
        RECT 213.675 58.145 213.935 58.405 ;
        RECT 213.675 57.485 213.935 57.745 ;
        RECT 213.675 56.825 213.935 57.085 ;
        RECT 213.675 56.165 213.935 56.425 ;
        RECT 213.675 55.505 213.935 55.765 ;
        RECT 213.675 54.845 213.935 55.105 ;
        RECT 213.675 54.185 213.935 54.445 ;
        RECT 213.675 53.525 213.935 53.785 ;
        RECT 213.675 52.865 213.935 53.125 ;
        RECT 213.675 52.205 213.935 52.465 ;
        RECT 213.675 51.545 213.935 51.805 ;
        RECT 213.675 50.885 213.935 51.145 ;
        RECT 213.675 50.225 213.935 50.485 ;
        RECT 218.160 47.865 218.420 48.125 ;
        RECT 218.820 47.865 219.080 48.125 ;
        RECT 219.480 47.865 219.740 48.125 ;
        RECT 218.160 47.205 218.420 47.465 ;
        RECT 218.820 47.205 219.080 47.465 ;
        RECT 219.480 47.205 219.740 47.465 ;
        RECT 218.160 46.545 218.420 46.805 ;
        RECT 218.820 46.545 219.080 46.805 ;
        RECT 219.480 46.545 219.740 46.805 ;
        RECT 218.160 22.265 218.420 22.525 ;
        RECT 218.820 22.265 219.080 22.525 ;
        RECT 219.480 22.265 219.740 22.525 ;
        RECT 218.160 21.605 218.420 21.865 ;
        RECT 218.820 21.605 219.080 21.865 ;
        RECT 219.480 21.605 219.740 21.865 ;
        RECT 218.160 20.945 218.420 21.205 ;
        RECT 218.820 20.945 219.080 21.205 ;
        RECT 219.480 20.945 219.740 21.205 ;
        RECT 223.965 58.805 224.225 59.065 ;
        RECT 223.965 58.145 224.225 58.405 ;
        RECT 223.965 57.485 224.225 57.745 ;
        RECT 223.965 56.825 224.225 57.085 ;
        RECT 223.965 56.165 224.225 56.425 ;
        RECT 223.965 55.505 224.225 55.765 ;
        RECT 223.965 54.845 224.225 55.105 ;
        RECT 223.965 54.185 224.225 54.445 ;
        RECT 223.965 53.525 224.225 53.785 ;
        RECT 223.965 52.865 224.225 53.125 ;
        RECT 223.965 52.205 224.225 52.465 ;
        RECT 223.965 51.545 224.225 51.805 ;
        RECT 223.965 50.885 224.225 51.145 ;
        RECT 223.965 50.225 224.225 50.485 ;
        RECT 235.615 59.990 235.875 60.250 ;
        RECT 253.460 59.990 253.720 60.250 ;
        RECT 228.460 45.165 228.720 45.425 ;
        RECT 229.120 45.165 229.380 45.425 ;
        RECT 229.780 45.165 230.040 45.425 ;
        RECT 228.460 44.505 228.720 44.765 ;
        RECT 229.120 44.505 229.380 44.765 ;
        RECT 229.780 44.505 230.040 44.765 ;
        RECT 228.460 43.845 228.720 44.105 ;
        RECT 229.120 43.845 229.380 44.105 ;
        RECT 229.780 43.845 230.040 44.105 ;
        RECT 228.460 24.965 228.720 25.225 ;
        RECT 229.120 24.965 229.380 25.225 ;
        RECT 229.780 24.965 230.040 25.225 ;
        RECT 228.460 24.305 228.720 24.565 ;
        RECT 229.120 24.305 229.380 24.565 ;
        RECT 229.780 24.305 230.040 24.565 ;
        RECT 228.460 23.645 228.720 23.905 ;
        RECT 229.120 23.645 229.380 23.905 ;
        RECT 229.780 23.645 230.040 23.905 ;
        RECT 203.335 8.805 203.595 9.065 ;
        RECT 222.600 8.805 222.860 9.065 ;
        RECT 234.250 58.805 234.510 59.065 ;
        RECT 234.250 58.145 234.510 58.405 ;
        RECT 234.250 57.485 234.510 57.745 ;
        RECT 234.250 56.825 234.510 57.085 ;
        RECT 234.250 56.165 234.510 56.425 ;
        RECT 234.250 55.505 234.510 55.765 ;
        RECT 234.250 54.845 234.510 55.105 ;
        RECT 234.250 54.185 234.510 54.445 ;
        RECT 234.250 53.525 234.510 53.785 ;
        RECT 234.250 52.865 234.510 53.125 ;
        RECT 234.250 52.205 234.510 52.465 ;
        RECT 234.250 51.545 234.510 51.805 ;
        RECT 234.250 50.885 234.510 51.145 ;
        RECT 234.250 50.225 234.510 50.485 ;
        RECT 238.735 42.465 238.995 42.725 ;
        RECT 239.395 42.465 239.655 42.725 ;
        RECT 240.055 42.465 240.315 42.725 ;
        RECT 238.735 41.805 238.995 42.065 ;
        RECT 239.395 41.805 239.655 42.065 ;
        RECT 240.055 41.805 240.315 42.065 ;
        RECT 238.735 41.145 238.995 41.405 ;
        RECT 239.395 41.145 239.655 41.405 ;
        RECT 240.055 41.145 240.315 41.405 ;
        RECT 238.735 27.665 238.995 27.925 ;
        RECT 239.395 27.665 239.655 27.925 ;
        RECT 240.055 27.665 240.315 27.925 ;
        RECT 238.735 27.005 238.995 27.265 ;
        RECT 239.395 27.005 239.655 27.265 ;
        RECT 240.055 27.005 240.315 27.265 ;
        RECT 238.735 26.345 238.995 26.605 ;
        RECT 239.395 26.345 239.655 26.605 ;
        RECT 240.055 26.345 240.315 26.605 ;
        RECT 244.540 58.805 244.800 59.065 ;
        RECT 244.540 58.145 244.800 58.405 ;
        RECT 244.540 57.485 244.800 57.745 ;
        RECT 244.540 56.825 244.800 57.085 ;
        RECT 244.540 56.165 244.800 56.425 ;
        RECT 244.540 55.505 244.800 55.765 ;
        RECT 244.540 54.845 244.800 55.105 ;
        RECT 244.540 54.185 244.800 54.445 ;
        RECT 244.540 53.525 244.800 53.785 ;
        RECT 244.540 52.865 244.800 53.125 ;
        RECT 244.540 52.205 244.800 52.465 ;
        RECT 244.540 51.545 244.800 51.805 ;
        RECT 244.540 50.885 244.800 51.145 ;
        RECT 244.540 50.225 244.800 50.485 ;
        RECT 257.610 59.990 257.870 60.250 ;
        RECT 275.455 59.990 275.715 60.250 ;
        RECT 249.035 39.765 249.295 40.025 ;
        RECT 249.695 39.765 249.955 40.025 ;
        RECT 250.355 39.765 250.615 40.025 ;
        RECT 249.035 39.105 249.295 39.365 ;
        RECT 249.695 39.105 249.955 39.365 ;
        RECT 250.355 39.105 250.615 39.365 ;
        RECT 249.035 38.445 249.295 38.705 ;
        RECT 249.695 38.445 249.955 38.705 ;
        RECT 250.355 38.445 250.615 38.705 ;
        RECT 249.035 30.365 249.295 30.625 ;
        RECT 249.695 30.365 249.955 30.625 ;
        RECT 250.355 30.365 250.615 30.625 ;
        RECT 249.035 29.705 249.295 29.965 ;
        RECT 249.695 29.705 249.955 29.965 ;
        RECT 250.355 29.705 250.615 29.965 ;
        RECT 249.035 29.045 249.295 29.305 ;
        RECT 249.695 29.045 249.955 29.305 ;
        RECT 250.355 29.045 250.615 29.305 ;
        RECT 225.330 8.805 225.590 9.065 ;
        RECT 243.175 8.805 243.435 9.065 ;
        RECT 254.825 58.805 255.085 59.065 ;
        RECT 254.825 58.145 255.085 58.405 ;
        RECT 254.825 57.485 255.085 57.745 ;
        RECT 254.825 56.825 255.085 57.085 ;
        RECT 254.825 56.165 255.085 56.425 ;
        RECT 254.825 55.505 255.085 55.765 ;
        RECT 254.825 54.845 255.085 55.105 ;
        RECT 254.825 54.185 255.085 54.445 ;
        RECT 254.825 53.525 255.085 53.785 ;
        RECT 254.825 52.865 255.085 53.125 ;
        RECT 254.825 52.205 255.085 52.465 ;
        RECT 254.825 51.545 255.085 51.805 ;
        RECT 254.825 50.885 255.085 51.145 ;
        RECT 254.825 50.225 255.085 50.485 ;
        RECT 256.245 58.805 256.505 59.065 ;
        RECT 256.245 58.145 256.505 58.405 ;
        RECT 256.245 57.485 256.505 57.745 ;
        RECT 256.245 56.825 256.505 57.085 ;
        RECT 256.245 56.165 256.505 56.425 ;
        RECT 256.245 55.505 256.505 55.765 ;
        RECT 256.245 54.845 256.505 55.105 ;
        RECT 256.245 54.185 256.505 54.445 ;
        RECT 256.245 53.525 256.505 53.785 ;
        RECT 256.245 52.865 256.505 53.125 ;
        RECT 256.245 52.205 256.505 52.465 ;
        RECT 256.245 51.545 256.505 51.805 ;
        RECT 256.245 50.885 256.505 51.145 ;
        RECT 256.245 50.225 256.505 50.485 ;
        RECT 260.730 47.865 260.990 48.125 ;
        RECT 261.390 47.865 261.650 48.125 ;
        RECT 262.050 47.865 262.310 48.125 ;
        RECT 260.730 47.205 260.990 47.465 ;
        RECT 261.390 47.205 261.650 47.465 ;
        RECT 262.050 47.205 262.310 47.465 ;
        RECT 260.730 46.545 260.990 46.805 ;
        RECT 261.390 46.545 261.650 46.805 ;
        RECT 262.050 46.545 262.310 46.805 ;
        RECT 260.730 22.265 260.990 22.525 ;
        RECT 261.390 22.265 261.650 22.525 ;
        RECT 262.050 22.265 262.310 22.525 ;
        RECT 260.730 21.605 260.990 21.865 ;
        RECT 261.390 21.605 261.650 21.865 ;
        RECT 262.050 21.605 262.310 21.865 ;
        RECT 260.730 20.945 260.990 21.205 ;
        RECT 261.390 20.945 261.650 21.205 ;
        RECT 262.050 20.945 262.310 21.205 ;
        RECT 266.535 58.805 266.795 59.065 ;
        RECT 266.535 58.145 266.795 58.405 ;
        RECT 266.535 57.485 266.795 57.745 ;
        RECT 266.535 56.825 266.795 57.085 ;
        RECT 266.535 56.165 266.795 56.425 ;
        RECT 266.535 55.505 266.795 55.765 ;
        RECT 266.535 54.845 266.795 55.105 ;
        RECT 266.535 54.185 266.795 54.445 ;
        RECT 266.535 53.525 266.795 53.785 ;
        RECT 266.535 52.865 266.795 53.125 ;
        RECT 266.535 52.205 266.795 52.465 ;
        RECT 266.535 51.545 266.795 51.805 ;
        RECT 266.535 50.885 266.795 51.145 ;
        RECT 266.535 50.225 266.795 50.485 ;
        RECT 278.185 59.990 278.445 60.250 ;
        RECT 296.030 59.990 296.290 60.250 ;
        RECT 271.030 45.165 271.290 45.425 ;
        RECT 271.690 45.165 271.950 45.425 ;
        RECT 272.350 45.165 272.610 45.425 ;
        RECT 271.030 44.505 271.290 44.765 ;
        RECT 271.690 44.505 271.950 44.765 ;
        RECT 272.350 44.505 272.610 44.765 ;
        RECT 271.030 43.845 271.290 44.105 ;
        RECT 271.690 43.845 271.950 44.105 ;
        RECT 272.350 43.845 272.610 44.105 ;
        RECT 271.030 24.965 271.290 25.225 ;
        RECT 271.690 24.965 271.950 25.225 ;
        RECT 272.350 24.965 272.610 25.225 ;
        RECT 271.030 24.305 271.290 24.565 ;
        RECT 271.690 24.305 271.950 24.565 ;
        RECT 272.350 24.305 272.610 24.565 ;
        RECT 271.030 23.645 271.290 23.905 ;
        RECT 271.690 23.645 271.950 23.905 ;
        RECT 272.350 23.645 272.610 23.905 ;
        RECT 245.905 8.805 246.165 9.065 ;
        RECT 265.170 8.805 265.430 9.065 ;
        RECT 276.820 58.805 277.080 59.065 ;
        RECT 276.820 58.145 277.080 58.405 ;
        RECT 276.820 57.485 277.080 57.745 ;
        RECT 276.820 56.825 277.080 57.085 ;
        RECT 276.820 56.165 277.080 56.425 ;
        RECT 276.820 55.505 277.080 55.765 ;
        RECT 276.820 54.845 277.080 55.105 ;
        RECT 276.820 54.185 277.080 54.445 ;
        RECT 276.820 53.525 277.080 53.785 ;
        RECT 276.820 52.865 277.080 53.125 ;
        RECT 276.820 52.205 277.080 52.465 ;
        RECT 276.820 51.545 277.080 51.805 ;
        RECT 276.820 50.885 277.080 51.145 ;
        RECT 276.820 50.225 277.080 50.485 ;
        RECT 281.305 42.465 281.565 42.725 ;
        RECT 281.965 42.465 282.225 42.725 ;
        RECT 282.625 42.465 282.885 42.725 ;
        RECT 281.305 41.805 281.565 42.065 ;
        RECT 281.965 41.805 282.225 42.065 ;
        RECT 282.625 41.805 282.885 42.065 ;
        RECT 281.305 41.145 281.565 41.405 ;
        RECT 281.965 41.145 282.225 41.405 ;
        RECT 282.625 41.145 282.885 41.405 ;
        RECT 281.305 27.665 281.565 27.925 ;
        RECT 281.965 27.665 282.225 27.925 ;
        RECT 282.625 27.665 282.885 27.925 ;
        RECT 281.305 27.005 281.565 27.265 ;
        RECT 281.965 27.005 282.225 27.265 ;
        RECT 282.625 27.005 282.885 27.265 ;
        RECT 281.305 26.345 281.565 26.605 ;
        RECT 281.965 26.345 282.225 26.605 ;
        RECT 282.625 26.345 282.885 26.605 ;
        RECT 287.110 58.805 287.370 59.065 ;
        RECT 287.110 58.145 287.370 58.405 ;
        RECT 287.110 57.485 287.370 57.745 ;
        RECT 287.110 56.825 287.370 57.085 ;
        RECT 287.110 56.165 287.370 56.425 ;
        RECT 287.110 55.505 287.370 55.765 ;
        RECT 287.110 54.845 287.370 55.105 ;
        RECT 287.110 54.185 287.370 54.445 ;
        RECT 287.110 53.525 287.370 53.785 ;
        RECT 287.110 52.865 287.370 53.125 ;
        RECT 287.110 52.205 287.370 52.465 ;
        RECT 287.110 51.545 287.370 51.805 ;
        RECT 287.110 50.885 287.370 51.145 ;
        RECT 287.110 50.225 287.370 50.485 ;
        RECT 300.180 59.990 300.440 60.250 ;
        RECT 318.025 59.990 318.285 60.250 ;
        RECT 291.605 39.765 291.865 40.025 ;
        RECT 292.265 39.765 292.525 40.025 ;
        RECT 292.925 39.765 293.185 40.025 ;
        RECT 291.605 39.105 291.865 39.365 ;
        RECT 292.265 39.105 292.525 39.365 ;
        RECT 292.925 39.105 293.185 39.365 ;
        RECT 291.605 38.445 291.865 38.705 ;
        RECT 292.265 38.445 292.525 38.705 ;
        RECT 292.925 38.445 293.185 38.705 ;
        RECT 291.605 30.365 291.865 30.625 ;
        RECT 292.265 30.365 292.525 30.625 ;
        RECT 292.925 30.365 293.185 30.625 ;
        RECT 291.605 29.705 291.865 29.965 ;
        RECT 292.265 29.705 292.525 29.965 ;
        RECT 292.925 29.705 293.185 29.965 ;
        RECT 291.605 29.045 291.865 29.305 ;
        RECT 292.265 29.045 292.525 29.305 ;
        RECT 292.925 29.045 293.185 29.305 ;
        RECT 267.900 8.805 268.160 9.065 ;
        RECT 285.745 8.805 286.005 9.065 ;
        RECT 297.395 58.805 297.655 59.065 ;
        RECT 297.395 58.145 297.655 58.405 ;
        RECT 297.395 57.485 297.655 57.745 ;
        RECT 297.395 56.825 297.655 57.085 ;
        RECT 297.395 56.165 297.655 56.425 ;
        RECT 297.395 55.505 297.655 55.765 ;
        RECT 297.395 54.845 297.655 55.105 ;
        RECT 297.395 54.185 297.655 54.445 ;
        RECT 297.395 53.525 297.655 53.785 ;
        RECT 297.395 52.865 297.655 53.125 ;
        RECT 297.395 52.205 297.655 52.465 ;
        RECT 297.395 51.545 297.655 51.805 ;
        RECT 297.395 50.885 297.655 51.145 ;
        RECT 297.395 50.225 297.655 50.485 ;
        RECT 298.815 58.805 299.075 59.065 ;
        RECT 298.815 58.145 299.075 58.405 ;
        RECT 298.815 57.485 299.075 57.745 ;
        RECT 298.815 56.825 299.075 57.085 ;
        RECT 298.815 56.165 299.075 56.425 ;
        RECT 298.815 55.505 299.075 55.765 ;
        RECT 298.815 54.845 299.075 55.105 ;
        RECT 298.815 54.185 299.075 54.445 ;
        RECT 298.815 53.525 299.075 53.785 ;
        RECT 298.815 52.865 299.075 53.125 ;
        RECT 298.815 52.205 299.075 52.465 ;
        RECT 298.815 51.545 299.075 51.805 ;
        RECT 298.815 50.885 299.075 51.145 ;
        RECT 298.815 50.225 299.075 50.485 ;
        RECT 303.300 47.865 303.560 48.125 ;
        RECT 303.960 47.865 304.220 48.125 ;
        RECT 304.620 47.865 304.880 48.125 ;
        RECT 303.300 47.205 303.560 47.465 ;
        RECT 303.960 47.205 304.220 47.465 ;
        RECT 304.620 47.205 304.880 47.465 ;
        RECT 303.300 46.545 303.560 46.805 ;
        RECT 303.960 46.545 304.220 46.805 ;
        RECT 304.620 46.545 304.880 46.805 ;
        RECT 303.300 22.265 303.560 22.525 ;
        RECT 303.960 22.265 304.220 22.525 ;
        RECT 304.620 22.265 304.880 22.525 ;
        RECT 303.300 21.605 303.560 21.865 ;
        RECT 303.960 21.605 304.220 21.865 ;
        RECT 304.620 21.605 304.880 21.865 ;
        RECT 303.300 20.945 303.560 21.205 ;
        RECT 303.960 20.945 304.220 21.205 ;
        RECT 304.620 20.945 304.880 21.205 ;
        RECT 309.105 58.805 309.365 59.065 ;
        RECT 309.105 58.145 309.365 58.405 ;
        RECT 309.105 57.485 309.365 57.745 ;
        RECT 309.105 56.825 309.365 57.085 ;
        RECT 309.105 56.165 309.365 56.425 ;
        RECT 309.105 55.505 309.365 55.765 ;
        RECT 309.105 54.845 309.365 55.105 ;
        RECT 309.105 54.185 309.365 54.445 ;
        RECT 309.105 53.525 309.365 53.785 ;
        RECT 309.105 52.865 309.365 53.125 ;
        RECT 309.105 52.205 309.365 52.465 ;
        RECT 309.105 51.545 309.365 51.805 ;
        RECT 309.105 50.885 309.365 51.145 ;
        RECT 309.105 50.225 309.365 50.485 ;
        RECT 320.755 59.990 321.015 60.250 ;
        RECT 338.600 59.990 338.860 60.250 ;
        RECT 313.600 45.165 313.860 45.425 ;
        RECT 314.260 45.165 314.520 45.425 ;
        RECT 314.920 45.165 315.180 45.425 ;
        RECT 313.600 44.505 313.860 44.765 ;
        RECT 314.260 44.505 314.520 44.765 ;
        RECT 314.920 44.505 315.180 44.765 ;
        RECT 313.600 43.845 313.860 44.105 ;
        RECT 314.260 43.845 314.520 44.105 ;
        RECT 314.920 43.845 315.180 44.105 ;
        RECT 313.600 24.965 313.860 25.225 ;
        RECT 314.260 24.965 314.520 25.225 ;
        RECT 314.920 24.965 315.180 25.225 ;
        RECT 313.600 24.305 313.860 24.565 ;
        RECT 314.260 24.305 314.520 24.565 ;
        RECT 314.920 24.305 315.180 24.565 ;
        RECT 313.600 23.645 313.860 23.905 ;
        RECT 314.260 23.645 314.520 23.905 ;
        RECT 314.920 23.645 315.180 23.905 ;
        RECT 288.475 8.805 288.735 9.065 ;
        RECT 307.740 8.805 308.000 9.065 ;
        RECT 319.390 58.805 319.650 59.065 ;
        RECT 319.390 58.145 319.650 58.405 ;
        RECT 319.390 57.485 319.650 57.745 ;
        RECT 319.390 56.825 319.650 57.085 ;
        RECT 319.390 56.165 319.650 56.425 ;
        RECT 319.390 55.505 319.650 55.765 ;
        RECT 319.390 54.845 319.650 55.105 ;
        RECT 319.390 54.185 319.650 54.445 ;
        RECT 319.390 53.525 319.650 53.785 ;
        RECT 319.390 52.865 319.650 53.125 ;
        RECT 319.390 52.205 319.650 52.465 ;
        RECT 319.390 51.545 319.650 51.805 ;
        RECT 319.390 50.885 319.650 51.145 ;
        RECT 319.390 50.225 319.650 50.485 ;
        RECT 323.875 42.465 324.135 42.725 ;
        RECT 324.535 42.465 324.795 42.725 ;
        RECT 325.195 42.465 325.455 42.725 ;
        RECT 323.875 41.805 324.135 42.065 ;
        RECT 324.535 41.805 324.795 42.065 ;
        RECT 325.195 41.805 325.455 42.065 ;
        RECT 323.875 41.145 324.135 41.405 ;
        RECT 324.535 41.145 324.795 41.405 ;
        RECT 325.195 41.145 325.455 41.405 ;
        RECT 323.875 27.665 324.135 27.925 ;
        RECT 324.535 27.665 324.795 27.925 ;
        RECT 325.195 27.665 325.455 27.925 ;
        RECT 323.875 27.005 324.135 27.265 ;
        RECT 324.535 27.005 324.795 27.265 ;
        RECT 325.195 27.005 325.455 27.265 ;
        RECT 323.875 26.345 324.135 26.605 ;
        RECT 324.535 26.345 324.795 26.605 ;
        RECT 325.195 26.345 325.455 26.605 ;
        RECT 329.680 58.805 329.940 59.065 ;
        RECT 329.680 58.145 329.940 58.405 ;
        RECT 329.680 57.485 329.940 57.745 ;
        RECT 329.680 56.825 329.940 57.085 ;
        RECT 329.680 56.165 329.940 56.425 ;
        RECT 329.680 55.505 329.940 55.765 ;
        RECT 329.680 54.845 329.940 55.105 ;
        RECT 329.680 54.185 329.940 54.445 ;
        RECT 329.680 53.525 329.940 53.785 ;
        RECT 329.680 52.865 329.940 53.125 ;
        RECT 329.680 52.205 329.940 52.465 ;
        RECT 329.680 51.545 329.940 51.805 ;
        RECT 329.680 50.885 329.940 51.145 ;
        RECT 329.680 50.225 329.940 50.485 ;
        RECT 342.750 59.990 343.010 60.250 ;
        RECT 360.595 59.990 360.855 60.250 ;
        RECT 334.175 39.765 334.435 40.025 ;
        RECT 334.835 39.765 335.095 40.025 ;
        RECT 335.495 39.765 335.755 40.025 ;
        RECT 334.175 39.105 334.435 39.365 ;
        RECT 334.835 39.105 335.095 39.365 ;
        RECT 335.495 39.105 335.755 39.365 ;
        RECT 334.175 38.445 334.435 38.705 ;
        RECT 334.835 38.445 335.095 38.705 ;
        RECT 335.495 38.445 335.755 38.705 ;
        RECT 334.175 30.365 334.435 30.625 ;
        RECT 334.835 30.365 335.095 30.625 ;
        RECT 335.495 30.365 335.755 30.625 ;
        RECT 334.175 29.705 334.435 29.965 ;
        RECT 334.835 29.705 335.095 29.965 ;
        RECT 335.495 29.705 335.755 29.965 ;
        RECT 334.175 29.045 334.435 29.305 ;
        RECT 334.835 29.045 335.095 29.305 ;
        RECT 335.495 29.045 335.755 29.305 ;
        RECT 310.470 8.805 310.730 9.065 ;
        RECT 328.315 8.805 328.575 9.065 ;
        RECT 339.965 58.805 340.225 59.065 ;
        RECT 339.965 58.145 340.225 58.405 ;
        RECT 339.965 57.485 340.225 57.745 ;
        RECT 339.965 56.825 340.225 57.085 ;
        RECT 339.965 56.165 340.225 56.425 ;
        RECT 339.965 55.505 340.225 55.765 ;
        RECT 339.965 54.845 340.225 55.105 ;
        RECT 339.965 54.185 340.225 54.445 ;
        RECT 339.965 53.525 340.225 53.785 ;
        RECT 339.965 52.865 340.225 53.125 ;
        RECT 339.965 52.205 340.225 52.465 ;
        RECT 339.965 51.545 340.225 51.805 ;
        RECT 339.965 50.885 340.225 51.145 ;
        RECT 339.965 50.225 340.225 50.485 ;
        RECT 341.385 58.805 341.645 59.065 ;
        RECT 341.385 58.145 341.645 58.405 ;
        RECT 341.385 57.485 341.645 57.745 ;
        RECT 341.385 56.825 341.645 57.085 ;
        RECT 341.385 56.165 341.645 56.425 ;
        RECT 341.385 55.505 341.645 55.765 ;
        RECT 341.385 54.845 341.645 55.105 ;
        RECT 341.385 54.185 341.645 54.445 ;
        RECT 341.385 53.525 341.645 53.785 ;
        RECT 341.385 52.865 341.645 53.125 ;
        RECT 341.385 52.205 341.645 52.465 ;
        RECT 341.385 51.545 341.645 51.805 ;
        RECT 341.385 50.885 341.645 51.145 ;
        RECT 341.385 50.225 341.645 50.485 ;
        RECT 345.870 47.865 346.130 48.125 ;
        RECT 346.530 47.865 346.790 48.125 ;
        RECT 347.190 47.865 347.450 48.125 ;
        RECT 345.870 47.205 346.130 47.465 ;
        RECT 346.530 47.205 346.790 47.465 ;
        RECT 347.190 47.205 347.450 47.465 ;
        RECT 345.870 46.545 346.130 46.805 ;
        RECT 346.530 46.545 346.790 46.805 ;
        RECT 347.190 46.545 347.450 46.805 ;
        RECT 345.870 22.265 346.130 22.525 ;
        RECT 346.530 22.265 346.790 22.525 ;
        RECT 347.190 22.265 347.450 22.525 ;
        RECT 345.870 21.605 346.130 21.865 ;
        RECT 346.530 21.605 346.790 21.865 ;
        RECT 347.190 21.605 347.450 21.865 ;
        RECT 345.870 20.945 346.130 21.205 ;
        RECT 346.530 20.945 346.790 21.205 ;
        RECT 347.190 20.945 347.450 21.205 ;
        RECT 351.675 58.805 351.935 59.065 ;
        RECT 351.675 58.145 351.935 58.405 ;
        RECT 351.675 57.485 351.935 57.745 ;
        RECT 351.675 56.825 351.935 57.085 ;
        RECT 351.675 56.165 351.935 56.425 ;
        RECT 351.675 55.505 351.935 55.765 ;
        RECT 351.675 54.845 351.935 55.105 ;
        RECT 351.675 54.185 351.935 54.445 ;
        RECT 351.675 53.525 351.935 53.785 ;
        RECT 351.675 52.865 351.935 53.125 ;
        RECT 351.675 52.205 351.935 52.465 ;
        RECT 351.675 51.545 351.935 51.805 ;
        RECT 351.675 50.885 351.935 51.145 ;
        RECT 351.675 50.225 351.935 50.485 ;
        RECT 363.325 59.990 363.585 60.250 ;
        RECT 381.170 59.990 381.430 60.250 ;
        RECT 356.170 45.165 356.430 45.425 ;
        RECT 356.830 45.165 357.090 45.425 ;
        RECT 357.490 45.165 357.750 45.425 ;
        RECT 356.170 44.505 356.430 44.765 ;
        RECT 356.830 44.505 357.090 44.765 ;
        RECT 357.490 44.505 357.750 44.765 ;
        RECT 356.170 43.845 356.430 44.105 ;
        RECT 356.830 43.845 357.090 44.105 ;
        RECT 357.490 43.845 357.750 44.105 ;
        RECT 356.170 24.965 356.430 25.225 ;
        RECT 356.830 24.965 357.090 25.225 ;
        RECT 357.490 24.965 357.750 25.225 ;
        RECT 356.170 24.305 356.430 24.565 ;
        RECT 356.830 24.305 357.090 24.565 ;
        RECT 357.490 24.305 357.750 24.565 ;
        RECT 356.170 23.645 356.430 23.905 ;
        RECT 356.830 23.645 357.090 23.905 ;
        RECT 357.490 23.645 357.750 23.905 ;
        RECT 331.045 8.805 331.305 9.065 ;
        RECT 350.310 8.805 350.570 9.065 ;
        RECT 361.960 58.805 362.220 59.065 ;
        RECT 361.960 58.145 362.220 58.405 ;
        RECT 361.960 57.485 362.220 57.745 ;
        RECT 361.960 56.825 362.220 57.085 ;
        RECT 361.960 56.165 362.220 56.425 ;
        RECT 361.960 55.505 362.220 55.765 ;
        RECT 361.960 54.845 362.220 55.105 ;
        RECT 361.960 54.185 362.220 54.445 ;
        RECT 361.960 53.525 362.220 53.785 ;
        RECT 361.960 52.865 362.220 53.125 ;
        RECT 361.960 52.205 362.220 52.465 ;
        RECT 361.960 51.545 362.220 51.805 ;
        RECT 361.960 50.885 362.220 51.145 ;
        RECT 361.960 50.225 362.220 50.485 ;
        RECT 366.445 42.465 366.705 42.725 ;
        RECT 367.105 42.465 367.365 42.725 ;
        RECT 367.765 42.465 368.025 42.725 ;
        RECT 366.445 41.805 366.705 42.065 ;
        RECT 367.105 41.805 367.365 42.065 ;
        RECT 367.765 41.805 368.025 42.065 ;
        RECT 366.445 41.145 366.705 41.405 ;
        RECT 367.105 41.145 367.365 41.405 ;
        RECT 367.765 41.145 368.025 41.405 ;
        RECT 366.445 27.665 366.705 27.925 ;
        RECT 367.105 27.665 367.365 27.925 ;
        RECT 367.765 27.665 368.025 27.925 ;
        RECT 366.445 27.005 366.705 27.265 ;
        RECT 367.105 27.005 367.365 27.265 ;
        RECT 367.765 27.005 368.025 27.265 ;
        RECT 366.445 26.345 366.705 26.605 ;
        RECT 367.105 26.345 367.365 26.605 ;
        RECT 367.765 26.345 368.025 26.605 ;
        RECT 372.250 58.805 372.510 59.065 ;
        RECT 372.250 58.145 372.510 58.405 ;
        RECT 372.250 57.485 372.510 57.745 ;
        RECT 372.250 56.825 372.510 57.085 ;
        RECT 372.250 56.165 372.510 56.425 ;
        RECT 372.250 55.505 372.510 55.765 ;
        RECT 372.250 54.845 372.510 55.105 ;
        RECT 372.250 54.185 372.510 54.445 ;
        RECT 372.250 53.525 372.510 53.785 ;
        RECT 372.250 52.865 372.510 53.125 ;
        RECT 372.250 52.205 372.510 52.465 ;
        RECT 372.250 51.545 372.510 51.805 ;
        RECT 372.250 50.885 372.510 51.145 ;
        RECT 372.250 50.225 372.510 50.485 ;
        RECT 385.320 59.990 385.580 60.250 ;
        RECT 403.165 59.990 403.425 60.250 ;
        RECT 376.745 39.765 377.005 40.025 ;
        RECT 377.405 39.765 377.665 40.025 ;
        RECT 378.065 39.765 378.325 40.025 ;
        RECT 376.745 39.105 377.005 39.365 ;
        RECT 377.405 39.105 377.665 39.365 ;
        RECT 378.065 39.105 378.325 39.365 ;
        RECT 376.745 38.445 377.005 38.705 ;
        RECT 377.405 38.445 377.665 38.705 ;
        RECT 378.065 38.445 378.325 38.705 ;
        RECT 376.745 30.365 377.005 30.625 ;
        RECT 377.405 30.365 377.665 30.625 ;
        RECT 378.065 30.365 378.325 30.625 ;
        RECT 376.745 29.705 377.005 29.965 ;
        RECT 377.405 29.705 377.665 29.965 ;
        RECT 378.065 29.705 378.325 29.965 ;
        RECT 376.745 29.045 377.005 29.305 ;
        RECT 377.405 29.045 377.665 29.305 ;
        RECT 378.065 29.045 378.325 29.305 ;
        RECT 353.040 8.805 353.300 9.065 ;
        RECT 370.885 8.805 371.145 9.065 ;
        RECT 382.535 58.805 382.795 59.065 ;
        RECT 382.535 58.145 382.795 58.405 ;
        RECT 382.535 57.485 382.795 57.745 ;
        RECT 382.535 56.825 382.795 57.085 ;
        RECT 382.535 56.165 382.795 56.425 ;
        RECT 382.535 55.505 382.795 55.765 ;
        RECT 382.535 54.845 382.795 55.105 ;
        RECT 382.535 54.185 382.795 54.445 ;
        RECT 382.535 53.525 382.795 53.785 ;
        RECT 382.535 52.865 382.795 53.125 ;
        RECT 382.535 52.205 382.795 52.465 ;
        RECT 382.535 51.545 382.795 51.805 ;
        RECT 382.535 50.885 382.795 51.145 ;
        RECT 382.535 50.225 382.795 50.485 ;
        RECT 383.955 58.805 384.215 59.065 ;
        RECT 383.955 58.145 384.215 58.405 ;
        RECT 383.955 57.485 384.215 57.745 ;
        RECT 383.955 56.825 384.215 57.085 ;
        RECT 383.955 56.165 384.215 56.425 ;
        RECT 383.955 55.505 384.215 55.765 ;
        RECT 383.955 54.845 384.215 55.105 ;
        RECT 383.955 54.185 384.215 54.445 ;
        RECT 383.955 53.525 384.215 53.785 ;
        RECT 383.955 52.865 384.215 53.125 ;
        RECT 383.955 52.205 384.215 52.465 ;
        RECT 383.955 51.545 384.215 51.805 ;
        RECT 383.955 50.885 384.215 51.145 ;
        RECT 383.955 50.225 384.215 50.485 ;
        RECT 388.440 47.865 388.700 48.125 ;
        RECT 389.100 47.865 389.360 48.125 ;
        RECT 389.760 47.865 390.020 48.125 ;
        RECT 388.440 47.205 388.700 47.465 ;
        RECT 389.100 47.205 389.360 47.465 ;
        RECT 389.760 47.205 390.020 47.465 ;
        RECT 388.440 46.545 388.700 46.805 ;
        RECT 389.100 46.545 389.360 46.805 ;
        RECT 389.760 46.545 390.020 46.805 ;
        RECT 388.440 22.265 388.700 22.525 ;
        RECT 389.100 22.265 389.360 22.525 ;
        RECT 389.760 22.265 390.020 22.525 ;
        RECT 388.440 21.605 388.700 21.865 ;
        RECT 389.100 21.605 389.360 21.865 ;
        RECT 389.760 21.605 390.020 21.865 ;
        RECT 388.440 20.945 388.700 21.205 ;
        RECT 389.100 20.945 389.360 21.205 ;
        RECT 389.760 20.945 390.020 21.205 ;
        RECT 394.245 58.805 394.505 59.065 ;
        RECT 394.245 58.145 394.505 58.405 ;
        RECT 394.245 57.485 394.505 57.745 ;
        RECT 394.245 56.825 394.505 57.085 ;
        RECT 394.245 56.165 394.505 56.425 ;
        RECT 394.245 55.505 394.505 55.765 ;
        RECT 394.245 54.845 394.505 55.105 ;
        RECT 394.245 54.185 394.505 54.445 ;
        RECT 394.245 53.525 394.505 53.785 ;
        RECT 394.245 52.865 394.505 53.125 ;
        RECT 394.245 52.205 394.505 52.465 ;
        RECT 394.245 51.545 394.505 51.805 ;
        RECT 394.245 50.885 394.505 51.145 ;
        RECT 394.245 50.225 394.505 50.485 ;
        RECT 405.895 59.990 406.155 60.250 ;
        RECT 423.740 59.990 424.000 60.250 ;
        RECT 398.740 45.165 399.000 45.425 ;
        RECT 399.400 45.165 399.660 45.425 ;
        RECT 400.060 45.165 400.320 45.425 ;
        RECT 398.740 44.505 399.000 44.765 ;
        RECT 399.400 44.505 399.660 44.765 ;
        RECT 400.060 44.505 400.320 44.765 ;
        RECT 398.740 43.845 399.000 44.105 ;
        RECT 399.400 43.845 399.660 44.105 ;
        RECT 400.060 43.845 400.320 44.105 ;
        RECT 398.740 24.965 399.000 25.225 ;
        RECT 399.400 24.965 399.660 25.225 ;
        RECT 400.060 24.965 400.320 25.225 ;
        RECT 398.740 24.305 399.000 24.565 ;
        RECT 399.400 24.305 399.660 24.565 ;
        RECT 400.060 24.305 400.320 24.565 ;
        RECT 398.740 23.645 399.000 23.905 ;
        RECT 399.400 23.645 399.660 23.905 ;
        RECT 400.060 23.645 400.320 23.905 ;
        RECT 373.615 8.805 373.875 9.065 ;
        RECT 392.880 8.805 393.140 9.065 ;
        RECT 404.530 58.805 404.790 59.065 ;
        RECT 404.530 58.145 404.790 58.405 ;
        RECT 404.530 57.485 404.790 57.745 ;
        RECT 404.530 56.825 404.790 57.085 ;
        RECT 404.530 56.165 404.790 56.425 ;
        RECT 404.530 55.505 404.790 55.765 ;
        RECT 404.530 54.845 404.790 55.105 ;
        RECT 404.530 54.185 404.790 54.445 ;
        RECT 404.530 53.525 404.790 53.785 ;
        RECT 404.530 52.865 404.790 53.125 ;
        RECT 404.530 52.205 404.790 52.465 ;
        RECT 404.530 51.545 404.790 51.805 ;
        RECT 404.530 50.885 404.790 51.145 ;
        RECT 404.530 50.225 404.790 50.485 ;
        RECT 409.015 42.465 409.275 42.725 ;
        RECT 409.675 42.465 409.935 42.725 ;
        RECT 410.335 42.465 410.595 42.725 ;
        RECT 409.015 41.805 409.275 42.065 ;
        RECT 409.675 41.805 409.935 42.065 ;
        RECT 410.335 41.805 410.595 42.065 ;
        RECT 409.015 41.145 409.275 41.405 ;
        RECT 409.675 41.145 409.935 41.405 ;
        RECT 410.335 41.145 410.595 41.405 ;
        RECT 409.015 27.665 409.275 27.925 ;
        RECT 409.675 27.665 409.935 27.925 ;
        RECT 410.335 27.665 410.595 27.925 ;
        RECT 409.015 27.005 409.275 27.265 ;
        RECT 409.675 27.005 409.935 27.265 ;
        RECT 410.335 27.005 410.595 27.265 ;
        RECT 409.015 26.345 409.275 26.605 ;
        RECT 409.675 26.345 409.935 26.605 ;
        RECT 410.335 26.345 410.595 26.605 ;
        RECT 414.820 58.805 415.080 59.065 ;
        RECT 414.820 58.145 415.080 58.405 ;
        RECT 414.820 57.485 415.080 57.745 ;
        RECT 414.820 56.825 415.080 57.085 ;
        RECT 414.820 56.165 415.080 56.425 ;
        RECT 414.820 55.505 415.080 55.765 ;
        RECT 414.820 54.845 415.080 55.105 ;
        RECT 414.820 54.185 415.080 54.445 ;
        RECT 414.820 53.525 415.080 53.785 ;
        RECT 414.820 52.865 415.080 53.125 ;
        RECT 414.820 52.205 415.080 52.465 ;
        RECT 414.820 51.545 415.080 51.805 ;
        RECT 414.820 50.885 415.080 51.145 ;
        RECT 414.820 50.225 415.080 50.485 ;
        RECT 427.890 59.990 428.150 60.250 ;
        RECT 445.735 59.990 445.995 60.250 ;
        RECT 419.315 39.765 419.575 40.025 ;
        RECT 419.975 39.765 420.235 40.025 ;
        RECT 420.635 39.765 420.895 40.025 ;
        RECT 419.315 39.105 419.575 39.365 ;
        RECT 419.975 39.105 420.235 39.365 ;
        RECT 420.635 39.105 420.895 39.365 ;
        RECT 419.315 38.445 419.575 38.705 ;
        RECT 419.975 38.445 420.235 38.705 ;
        RECT 420.635 38.445 420.895 38.705 ;
        RECT 419.315 30.365 419.575 30.625 ;
        RECT 419.975 30.365 420.235 30.625 ;
        RECT 420.635 30.365 420.895 30.625 ;
        RECT 419.315 29.705 419.575 29.965 ;
        RECT 419.975 29.705 420.235 29.965 ;
        RECT 420.635 29.705 420.895 29.965 ;
        RECT 419.315 29.045 419.575 29.305 ;
        RECT 419.975 29.045 420.235 29.305 ;
        RECT 420.635 29.045 420.895 29.305 ;
        RECT 395.610 8.805 395.870 9.065 ;
        RECT 413.455 8.805 413.715 9.065 ;
        RECT 425.105 58.805 425.365 59.065 ;
        RECT 425.105 58.145 425.365 58.405 ;
        RECT 425.105 57.485 425.365 57.745 ;
        RECT 425.105 56.825 425.365 57.085 ;
        RECT 425.105 56.165 425.365 56.425 ;
        RECT 425.105 55.505 425.365 55.765 ;
        RECT 425.105 54.845 425.365 55.105 ;
        RECT 425.105 54.185 425.365 54.445 ;
        RECT 425.105 53.525 425.365 53.785 ;
        RECT 425.105 52.865 425.365 53.125 ;
        RECT 425.105 52.205 425.365 52.465 ;
        RECT 425.105 51.545 425.365 51.805 ;
        RECT 425.105 50.885 425.365 51.145 ;
        RECT 425.105 50.225 425.365 50.485 ;
        RECT 426.525 58.805 426.785 59.065 ;
        RECT 426.525 58.145 426.785 58.405 ;
        RECT 426.525 57.485 426.785 57.745 ;
        RECT 426.525 56.825 426.785 57.085 ;
        RECT 426.525 56.165 426.785 56.425 ;
        RECT 426.525 55.505 426.785 55.765 ;
        RECT 426.525 54.845 426.785 55.105 ;
        RECT 426.525 54.185 426.785 54.445 ;
        RECT 426.525 53.525 426.785 53.785 ;
        RECT 426.525 52.865 426.785 53.125 ;
        RECT 426.525 52.205 426.785 52.465 ;
        RECT 426.525 51.545 426.785 51.805 ;
        RECT 426.525 50.885 426.785 51.145 ;
        RECT 426.525 50.225 426.785 50.485 ;
        RECT 431.010 47.865 431.270 48.125 ;
        RECT 431.670 47.865 431.930 48.125 ;
        RECT 432.330 47.865 432.590 48.125 ;
        RECT 431.010 47.205 431.270 47.465 ;
        RECT 431.670 47.205 431.930 47.465 ;
        RECT 432.330 47.205 432.590 47.465 ;
        RECT 431.010 46.545 431.270 46.805 ;
        RECT 431.670 46.545 431.930 46.805 ;
        RECT 432.330 46.545 432.590 46.805 ;
        RECT 431.010 22.265 431.270 22.525 ;
        RECT 431.670 22.265 431.930 22.525 ;
        RECT 432.330 22.265 432.590 22.525 ;
        RECT 431.010 21.605 431.270 21.865 ;
        RECT 431.670 21.605 431.930 21.865 ;
        RECT 432.330 21.605 432.590 21.865 ;
        RECT 431.010 20.945 431.270 21.205 ;
        RECT 431.670 20.945 431.930 21.205 ;
        RECT 432.330 20.945 432.590 21.205 ;
        RECT 436.815 58.805 437.075 59.065 ;
        RECT 436.815 58.145 437.075 58.405 ;
        RECT 436.815 57.485 437.075 57.745 ;
        RECT 436.815 56.825 437.075 57.085 ;
        RECT 436.815 56.165 437.075 56.425 ;
        RECT 436.815 55.505 437.075 55.765 ;
        RECT 436.815 54.845 437.075 55.105 ;
        RECT 436.815 54.185 437.075 54.445 ;
        RECT 436.815 53.525 437.075 53.785 ;
        RECT 436.815 52.865 437.075 53.125 ;
        RECT 436.815 52.205 437.075 52.465 ;
        RECT 436.815 51.545 437.075 51.805 ;
        RECT 436.815 50.885 437.075 51.145 ;
        RECT 436.815 50.225 437.075 50.485 ;
        RECT 448.465 59.990 448.725 60.250 ;
        RECT 466.310 59.990 466.570 60.250 ;
        RECT 441.310 45.165 441.570 45.425 ;
        RECT 441.970 45.165 442.230 45.425 ;
        RECT 442.630 45.165 442.890 45.425 ;
        RECT 441.310 44.505 441.570 44.765 ;
        RECT 441.970 44.505 442.230 44.765 ;
        RECT 442.630 44.505 442.890 44.765 ;
        RECT 441.310 43.845 441.570 44.105 ;
        RECT 441.970 43.845 442.230 44.105 ;
        RECT 442.630 43.845 442.890 44.105 ;
        RECT 441.310 24.965 441.570 25.225 ;
        RECT 441.970 24.965 442.230 25.225 ;
        RECT 442.630 24.965 442.890 25.225 ;
        RECT 441.310 24.305 441.570 24.565 ;
        RECT 441.970 24.305 442.230 24.565 ;
        RECT 442.630 24.305 442.890 24.565 ;
        RECT 441.310 23.645 441.570 23.905 ;
        RECT 441.970 23.645 442.230 23.905 ;
        RECT 442.630 23.645 442.890 23.905 ;
        RECT 416.185 8.805 416.445 9.065 ;
        RECT 435.450 8.805 435.710 9.065 ;
        RECT 447.100 58.805 447.360 59.065 ;
        RECT 447.100 58.145 447.360 58.405 ;
        RECT 447.100 57.485 447.360 57.745 ;
        RECT 447.100 56.825 447.360 57.085 ;
        RECT 447.100 56.165 447.360 56.425 ;
        RECT 447.100 55.505 447.360 55.765 ;
        RECT 447.100 54.845 447.360 55.105 ;
        RECT 447.100 54.185 447.360 54.445 ;
        RECT 447.100 53.525 447.360 53.785 ;
        RECT 447.100 52.865 447.360 53.125 ;
        RECT 447.100 52.205 447.360 52.465 ;
        RECT 447.100 51.545 447.360 51.805 ;
        RECT 447.100 50.885 447.360 51.145 ;
        RECT 447.100 50.225 447.360 50.485 ;
        RECT 451.585 42.465 451.845 42.725 ;
        RECT 452.245 42.465 452.505 42.725 ;
        RECT 452.905 42.465 453.165 42.725 ;
        RECT 451.585 41.805 451.845 42.065 ;
        RECT 452.245 41.805 452.505 42.065 ;
        RECT 452.905 41.805 453.165 42.065 ;
        RECT 451.585 41.145 451.845 41.405 ;
        RECT 452.245 41.145 452.505 41.405 ;
        RECT 452.905 41.145 453.165 41.405 ;
        RECT 451.585 27.665 451.845 27.925 ;
        RECT 452.245 27.665 452.505 27.925 ;
        RECT 452.905 27.665 453.165 27.925 ;
        RECT 451.585 27.005 451.845 27.265 ;
        RECT 452.245 27.005 452.505 27.265 ;
        RECT 452.905 27.005 453.165 27.265 ;
        RECT 451.585 26.345 451.845 26.605 ;
        RECT 452.245 26.345 452.505 26.605 ;
        RECT 452.905 26.345 453.165 26.605 ;
        RECT 457.390 58.805 457.650 59.065 ;
        RECT 457.390 58.145 457.650 58.405 ;
        RECT 457.390 57.485 457.650 57.745 ;
        RECT 457.390 56.825 457.650 57.085 ;
        RECT 457.390 56.165 457.650 56.425 ;
        RECT 457.390 55.505 457.650 55.765 ;
        RECT 457.390 54.845 457.650 55.105 ;
        RECT 457.390 54.185 457.650 54.445 ;
        RECT 457.390 53.525 457.650 53.785 ;
        RECT 457.390 52.865 457.650 53.125 ;
        RECT 457.390 52.205 457.650 52.465 ;
        RECT 457.390 51.545 457.650 51.805 ;
        RECT 457.390 50.885 457.650 51.145 ;
        RECT 457.390 50.225 457.650 50.485 ;
        RECT 470.460 59.990 470.720 60.250 ;
        RECT 488.305 59.990 488.565 60.250 ;
        RECT 461.885 39.765 462.145 40.025 ;
        RECT 462.545 39.765 462.805 40.025 ;
        RECT 463.205 39.765 463.465 40.025 ;
        RECT 461.885 39.105 462.145 39.365 ;
        RECT 462.545 39.105 462.805 39.365 ;
        RECT 463.205 39.105 463.465 39.365 ;
        RECT 461.885 38.445 462.145 38.705 ;
        RECT 462.545 38.445 462.805 38.705 ;
        RECT 463.205 38.445 463.465 38.705 ;
        RECT 461.885 30.365 462.145 30.625 ;
        RECT 462.545 30.365 462.805 30.625 ;
        RECT 463.205 30.365 463.465 30.625 ;
        RECT 461.885 29.705 462.145 29.965 ;
        RECT 462.545 29.705 462.805 29.965 ;
        RECT 463.205 29.705 463.465 29.965 ;
        RECT 461.885 29.045 462.145 29.305 ;
        RECT 462.545 29.045 462.805 29.305 ;
        RECT 463.205 29.045 463.465 29.305 ;
        RECT 438.180 8.805 438.440 9.065 ;
        RECT 456.025 8.805 456.285 9.065 ;
        RECT 467.675 58.805 467.935 59.065 ;
        RECT 467.675 58.145 467.935 58.405 ;
        RECT 467.675 57.485 467.935 57.745 ;
        RECT 467.675 56.825 467.935 57.085 ;
        RECT 467.675 56.165 467.935 56.425 ;
        RECT 467.675 55.505 467.935 55.765 ;
        RECT 467.675 54.845 467.935 55.105 ;
        RECT 467.675 54.185 467.935 54.445 ;
        RECT 467.675 53.525 467.935 53.785 ;
        RECT 467.675 52.865 467.935 53.125 ;
        RECT 467.675 52.205 467.935 52.465 ;
        RECT 467.675 51.545 467.935 51.805 ;
        RECT 467.675 50.885 467.935 51.145 ;
        RECT 467.675 50.225 467.935 50.485 ;
        RECT 469.095 58.805 469.355 59.065 ;
        RECT 469.095 58.145 469.355 58.405 ;
        RECT 469.095 57.485 469.355 57.745 ;
        RECT 469.095 56.825 469.355 57.085 ;
        RECT 469.095 56.165 469.355 56.425 ;
        RECT 469.095 55.505 469.355 55.765 ;
        RECT 469.095 54.845 469.355 55.105 ;
        RECT 469.095 54.185 469.355 54.445 ;
        RECT 469.095 53.525 469.355 53.785 ;
        RECT 469.095 52.865 469.355 53.125 ;
        RECT 469.095 52.205 469.355 52.465 ;
        RECT 469.095 51.545 469.355 51.805 ;
        RECT 469.095 50.885 469.355 51.145 ;
        RECT 469.095 50.225 469.355 50.485 ;
        RECT 473.580 47.865 473.840 48.125 ;
        RECT 474.240 47.865 474.500 48.125 ;
        RECT 474.900 47.865 475.160 48.125 ;
        RECT 473.580 47.205 473.840 47.465 ;
        RECT 474.240 47.205 474.500 47.465 ;
        RECT 474.900 47.205 475.160 47.465 ;
        RECT 473.580 46.545 473.840 46.805 ;
        RECT 474.240 46.545 474.500 46.805 ;
        RECT 474.900 46.545 475.160 46.805 ;
        RECT 473.580 22.265 473.840 22.525 ;
        RECT 474.240 22.265 474.500 22.525 ;
        RECT 474.900 22.265 475.160 22.525 ;
        RECT 473.580 21.605 473.840 21.865 ;
        RECT 474.240 21.605 474.500 21.865 ;
        RECT 474.900 21.605 475.160 21.865 ;
        RECT 473.580 20.945 473.840 21.205 ;
        RECT 474.240 20.945 474.500 21.205 ;
        RECT 474.900 20.945 475.160 21.205 ;
        RECT 479.385 58.805 479.645 59.065 ;
        RECT 479.385 58.145 479.645 58.405 ;
        RECT 479.385 57.485 479.645 57.745 ;
        RECT 479.385 56.825 479.645 57.085 ;
        RECT 479.385 56.165 479.645 56.425 ;
        RECT 479.385 55.505 479.645 55.765 ;
        RECT 479.385 54.845 479.645 55.105 ;
        RECT 479.385 54.185 479.645 54.445 ;
        RECT 479.385 53.525 479.645 53.785 ;
        RECT 479.385 52.865 479.645 53.125 ;
        RECT 479.385 52.205 479.645 52.465 ;
        RECT 479.385 51.545 479.645 51.805 ;
        RECT 479.385 50.885 479.645 51.145 ;
        RECT 479.385 50.225 479.645 50.485 ;
        RECT 491.035 59.990 491.295 60.250 ;
        RECT 508.880 59.990 509.140 60.250 ;
        RECT 483.880 45.165 484.140 45.425 ;
        RECT 484.540 45.165 484.800 45.425 ;
        RECT 485.200 45.165 485.460 45.425 ;
        RECT 483.880 44.505 484.140 44.765 ;
        RECT 484.540 44.505 484.800 44.765 ;
        RECT 485.200 44.505 485.460 44.765 ;
        RECT 483.880 43.845 484.140 44.105 ;
        RECT 484.540 43.845 484.800 44.105 ;
        RECT 485.200 43.845 485.460 44.105 ;
        RECT 483.880 24.965 484.140 25.225 ;
        RECT 484.540 24.965 484.800 25.225 ;
        RECT 485.200 24.965 485.460 25.225 ;
        RECT 483.880 24.305 484.140 24.565 ;
        RECT 484.540 24.305 484.800 24.565 ;
        RECT 485.200 24.305 485.460 24.565 ;
        RECT 483.880 23.645 484.140 23.905 ;
        RECT 484.540 23.645 484.800 23.905 ;
        RECT 485.200 23.645 485.460 23.905 ;
        RECT 458.755 8.805 459.015 9.065 ;
        RECT 478.020 8.805 478.280 9.065 ;
        RECT 489.670 58.805 489.930 59.065 ;
        RECT 489.670 58.145 489.930 58.405 ;
        RECT 489.670 57.485 489.930 57.745 ;
        RECT 489.670 56.825 489.930 57.085 ;
        RECT 489.670 56.165 489.930 56.425 ;
        RECT 489.670 55.505 489.930 55.765 ;
        RECT 489.670 54.845 489.930 55.105 ;
        RECT 489.670 54.185 489.930 54.445 ;
        RECT 489.670 53.525 489.930 53.785 ;
        RECT 489.670 52.865 489.930 53.125 ;
        RECT 489.670 52.205 489.930 52.465 ;
        RECT 489.670 51.545 489.930 51.805 ;
        RECT 489.670 50.885 489.930 51.145 ;
        RECT 489.670 50.225 489.930 50.485 ;
        RECT 494.155 42.465 494.415 42.725 ;
        RECT 494.815 42.465 495.075 42.725 ;
        RECT 495.475 42.465 495.735 42.725 ;
        RECT 494.155 41.805 494.415 42.065 ;
        RECT 494.815 41.805 495.075 42.065 ;
        RECT 495.475 41.805 495.735 42.065 ;
        RECT 494.155 41.145 494.415 41.405 ;
        RECT 494.815 41.145 495.075 41.405 ;
        RECT 495.475 41.145 495.735 41.405 ;
        RECT 494.155 27.665 494.415 27.925 ;
        RECT 494.815 27.665 495.075 27.925 ;
        RECT 495.475 27.665 495.735 27.925 ;
        RECT 494.155 27.005 494.415 27.265 ;
        RECT 494.815 27.005 495.075 27.265 ;
        RECT 495.475 27.005 495.735 27.265 ;
        RECT 494.155 26.345 494.415 26.605 ;
        RECT 494.815 26.345 495.075 26.605 ;
        RECT 495.475 26.345 495.735 26.605 ;
        RECT 499.960 58.805 500.220 59.065 ;
        RECT 499.960 58.145 500.220 58.405 ;
        RECT 499.960 57.485 500.220 57.745 ;
        RECT 499.960 56.825 500.220 57.085 ;
        RECT 499.960 56.165 500.220 56.425 ;
        RECT 499.960 55.505 500.220 55.765 ;
        RECT 499.960 54.845 500.220 55.105 ;
        RECT 499.960 54.185 500.220 54.445 ;
        RECT 499.960 53.525 500.220 53.785 ;
        RECT 499.960 52.865 500.220 53.125 ;
        RECT 499.960 52.205 500.220 52.465 ;
        RECT 499.960 51.545 500.220 51.805 ;
        RECT 499.960 50.885 500.220 51.145 ;
        RECT 499.960 50.225 500.220 50.485 ;
        RECT 513.030 59.990 513.290 60.250 ;
        RECT 530.875 59.990 531.135 60.250 ;
        RECT 504.455 39.765 504.715 40.025 ;
        RECT 505.115 39.765 505.375 40.025 ;
        RECT 505.775 39.765 506.035 40.025 ;
        RECT 504.455 39.105 504.715 39.365 ;
        RECT 505.115 39.105 505.375 39.365 ;
        RECT 505.775 39.105 506.035 39.365 ;
        RECT 504.455 38.445 504.715 38.705 ;
        RECT 505.115 38.445 505.375 38.705 ;
        RECT 505.775 38.445 506.035 38.705 ;
        RECT 504.455 30.365 504.715 30.625 ;
        RECT 505.115 30.365 505.375 30.625 ;
        RECT 505.775 30.365 506.035 30.625 ;
        RECT 504.455 29.705 504.715 29.965 ;
        RECT 505.115 29.705 505.375 29.965 ;
        RECT 505.775 29.705 506.035 29.965 ;
        RECT 504.455 29.045 504.715 29.305 ;
        RECT 505.115 29.045 505.375 29.305 ;
        RECT 505.775 29.045 506.035 29.305 ;
        RECT 480.750 8.805 481.010 9.065 ;
        RECT 498.595 8.805 498.855 9.065 ;
        RECT 510.245 58.805 510.505 59.065 ;
        RECT 510.245 58.145 510.505 58.405 ;
        RECT 510.245 57.485 510.505 57.745 ;
        RECT 510.245 56.825 510.505 57.085 ;
        RECT 510.245 56.165 510.505 56.425 ;
        RECT 510.245 55.505 510.505 55.765 ;
        RECT 510.245 54.845 510.505 55.105 ;
        RECT 510.245 54.185 510.505 54.445 ;
        RECT 510.245 53.525 510.505 53.785 ;
        RECT 510.245 52.865 510.505 53.125 ;
        RECT 510.245 52.205 510.505 52.465 ;
        RECT 510.245 51.545 510.505 51.805 ;
        RECT 510.245 50.885 510.505 51.145 ;
        RECT 510.245 50.225 510.505 50.485 ;
        RECT 511.665 58.805 511.925 59.065 ;
        RECT 511.665 58.145 511.925 58.405 ;
        RECT 511.665 57.485 511.925 57.745 ;
        RECT 511.665 56.825 511.925 57.085 ;
        RECT 511.665 56.165 511.925 56.425 ;
        RECT 511.665 55.505 511.925 55.765 ;
        RECT 511.665 54.845 511.925 55.105 ;
        RECT 511.665 54.185 511.925 54.445 ;
        RECT 511.665 53.525 511.925 53.785 ;
        RECT 511.665 52.865 511.925 53.125 ;
        RECT 511.665 52.205 511.925 52.465 ;
        RECT 511.665 51.545 511.925 51.805 ;
        RECT 511.665 50.885 511.925 51.145 ;
        RECT 511.665 50.225 511.925 50.485 ;
        RECT 516.150 47.865 516.410 48.125 ;
        RECT 516.810 47.865 517.070 48.125 ;
        RECT 517.470 47.865 517.730 48.125 ;
        RECT 516.150 47.205 516.410 47.465 ;
        RECT 516.810 47.205 517.070 47.465 ;
        RECT 517.470 47.205 517.730 47.465 ;
        RECT 516.150 46.545 516.410 46.805 ;
        RECT 516.810 46.545 517.070 46.805 ;
        RECT 517.470 46.545 517.730 46.805 ;
        RECT 516.150 22.265 516.410 22.525 ;
        RECT 516.810 22.265 517.070 22.525 ;
        RECT 517.470 22.265 517.730 22.525 ;
        RECT 516.150 21.605 516.410 21.865 ;
        RECT 516.810 21.605 517.070 21.865 ;
        RECT 517.470 21.605 517.730 21.865 ;
        RECT 516.150 20.945 516.410 21.205 ;
        RECT 516.810 20.945 517.070 21.205 ;
        RECT 517.470 20.945 517.730 21.205 ;
        RECT 521.955 58.805 522.215 59.065 ;
        RECT 521.955 58.145 522.215 58.405 ;
        RECT 521.955 57.485 522.215 57.745 ;
        RECT 521.955 56.825 522.215 57.085 ;
        RECT 521.955 56.165 522.215 56.425 ;
        RECT 521.955 55.505 522.215 55.765 ;
        RECT 521.955 54.845 522.215 55.105 ;
        RECT 521.955 54.185 522.215 54.445 ;
        RECT 521.955 53.525 522.215 53.785 ;
        RECT 521.955 52.865 522.215 53.125 ;
        RECT 521.955 52.205 522.215 52.465 ;
        RECT 521.955 51.545 522.215 51.805 ;
        RECT 521.955 50.885 522.215 51.145 ;
        RECT 521.955 50.225 522.215 50.485 ;
        RECT 533.605 59.990 533.865 60.250 ;
        RECT 551.450 59.990 551.710 60.250 ;
        RECT 526.450 45.165 526.710 45.425 ;
        RECT 527.110 45.165 527.370 45.425 ;
        RECT 527.770 45.165 528.030 45.425 ;
        RECT 526.450 44.505 526.710 44.765 ;
        RECT 527.110 44.505 527.370 44.765 ;
        RECT 527.770 44.505 528.030 44.765 ;
        RECT 526.450 43.845 526.710 44.105 ;
        RECT 527.110 43.845 527.370 44.105 ;
        RECT 527.770 43.845 528.030 44.105 ;
        RECT 526.450 24.965 526.710 25.225 ;
        RECT 527.110 24.965 527.370 25.225 ;
        RECT 527.770 24.965 528.030 25.225 ;
        RECT 526.450 24.305 526.710 24.565 ;
        RECT 527.110 24.305 527.370 24.565 ;
        RECT 527.770 24.305 528.030 24.565 ;
        RECT 526.450 23.645 526.710 23.905 ;
        RECT 527.110 23.645 527.370 23.905 ;
        RECT 527.770 23.645 528.030 23.905 ;
        RECT 501.325 8.805 501.585 9.065 ;
        RECT 520.590 8.805 520.850 9.065 ;
        RECT 532.240 58.805 532.500 59.065 ;
        RECT 532.240 58.145 532.500 58.405 ;
        RECT 532.240 57.485 532.500 57.745 ;
        RECT 532.240 56.825 532.500 57.085 ;
        RECT 532.240 56.165 532.500 56.425 ;
        RECT 532.240 55.505 532.500 55.765 ;
        RECT 532.240 54.845 532.500 55.105 ;
        RECT 532.240 54.185 532.500 54.445 ;
        RECT 532.240 53.525 532.500 53.785 ;
        RECT 532.240 52.865 532.500 53.125 ;
        RECT 532.240 52.205 532.500 52.465 ;
        RECT 532.240 51.545 532.500 51.805 ;
        RECT 532.240 50.885 532.500 51.145 ;
        RECT 532.240 50.225 532.500 50.485 ;
        RECT 536.725 42.465 536.985 42.725 ;
        RECT 537.385 42.465 537.645 42.725 ;
        RECT 538.045 42.465 538.305 42.725 ;
        RECT 536.725 41.805 536.985 42.065 ;
        RECT 537.385 41.805 537.645 42.065 ;
        RECT 538.045 41.805 538.305 42.065 ;
        RECT 536.725 41.145 536.985 41.405 ;
        RECT 537.385 41.145 537.645 41.405 ;
        RECT 538.045 41.145 538.305 41.405 ;
        RECT 536.725 27.665 536.985 27.925 ;
        RECT 537.385 27.665 537.645 27.925 ;
        RECT 538.045 27.665 538.305 27.925 ;
        RECT 536.725 27.005 536.985 27.265 ;
        RECT 537.385 27.005 537.645 27.265 ;
        RECT 538.045 27.005 538.305 27.265 ;
        RECT 536.725 26.345 536.985 26.605 ;
        RECT 537.385 26.345 537.645 26.605 ;
        RECT 538.045 26.345 538.305 26.605 ;
        RECT 542.530 58.805 542.790 59.065 ;
        RECT 542.530 58.145 542.790 58.405 ;
        RECT 542.530 57.485 542.790 57.745 ;
        RECT 542.530 56.825 542.790 57.085 ;
        RECT 542.530 56.165 542.790 56.425 ;
        RECT 542.530 55.505 542.790 55.765 ;
        RECT 542.530 54.845 542.790 55.105 ;
        RECT 542.530 54.185 542.790 54.445 ;
        RECT 542.530 53.525 542.790 53.785 ;
        RECT 542.530 52.865 542.790 53.125 ;
        RECT 542.530 52.205 542.790 52.465 ;
        RECT 542.530 51.545 542.790 51.805 ;
        RECT 542.530 50.885 542.790 51.145 ;
        RECT 542.530 50.225 542.790 50.485 ;
        RECT 555.600 59.990 555.860 60.250 ;
        RECT 573.445 59.990 573.705 60.250 ;
        RECT 547.025 39.765 547.285 40.025 ;
        RECT 547.685 39.765 547.945 40.025 ;
        RECT 548.345 39.765 548.605 40.025 ;
        RECT 547.025 39.105 547.285 39.365 ;
        RECT 547.685 39.105 547.945 39.365 ;
        RECT 548.345 39.105 548.605 39.365 ;
        RECT 547.025 38.445 547.285 38.705 ;
        RECT 547.685 38.445 547.945 38.705 ;
        RECT 548.345 38.445 548.605 38.705 ;
        RECT 547.025 30.365 547.285 30.625 ;
        RECT 547.685 30.365 547.945 30.625 ;
        RECT 548.345 30.365 548.605 30.625 ;
        RECT 547.025 29.705 547.285 29.965 ;
        RECT 547.685 29.705 547.945 29.965 ;
        RECT 548.345 29.705 548.605 29.965 ;
        RECT 547.025 29.045 547.285 29.305 ;
        RECT 547.685 29.045 547.945 29.305 ;
        RECT 548.345 29.045 548.605 29.305 ;
        RECT 523.320 8.805 523.580 9.065 ;
        RECT 541.165 8.805 541.425 9.065 ;
        RECT 552.815 58.805 553.075 59.065 ;
        RECT 552.815 58.145 553.075 58.405 ;
        RECT 552.815 57.485 553.075 57.745 ;
        RECT 552.815 56.825 553.075 57.085 ;
        RECT 552.815 56.165 553.075 56.425 ;
        RECT 552.815 55.505 553.075 55.765 ;
        RECT 552.815 54.845 553.075 55.105 ;
        RECT 552.815 54.185 553.075 54.445 ;
        RECT 552.815 53.525 553.075 53.785 ;
        RECT 552.815 52.865 553.075 53.125 ;
        RECT 552.815 52.205 553.075 52.465 ;
        RECT 552.815 51.545 553.075 51.805 ;
        RECT 552.815 50.885 553.075 51.145 ;
        RECT 552.815 50.225 553.075 50.485 ;
        RECT 554.235 58.805 554.495 59.065 ;
        RECT 554.235 58.145 554.495 58.405 ;
        RECT 554.235 57.485 554.495 57.745 ;
        RECT 554.235 56.825 554.495 57.085 ;
        RECT 554.235 56.165 554.495 56.425 ;
        RECT 554.235 55.505 554.495 55.765 ;
        RECT 554.235 54.845 554.495 55.105 ;
        RECT 554.235 54.185 554.495 54.445 ;
        RECT 554.235 53.525 554.495 53.785 ;
        RECT 554.235 52.865 554.495 53.125 ;
        RECT 554.235 52.205 554.495 52.465 ;
        RECT 554.235 51.545 554.495 51.805 ;
        RECT 554.235 50.885 554.495 51.145 ;
        RECT 554.235 50.225 554.495 50.485 ;
        RECT 558.720 47.865 558.980 48.125 ;
        RECT 559.380 47.865 559.640 48.125 ;
        RECT 560.040 47.865 560.300 48.125 ;
        RECT 558.720 47.205 558.980 47.465 ;
        RECT 559.380 47.205 559.640 47.465 ;
        RECT 560.040 47.205 560.300 47.465 ;
        RECT 558.720 46.545 558.980 46.805 ;
        RECT 559.380 46.545 559.640 46.805 ;
        RECT 560.040 46.545 560.300 46.805 ;
        RECT 558.720 22.265 558.980 22.525 ;
        RECT 559.380 22.265 559.640 22.525 ;
        RECT 560.040 22.265 560.300 22.525 ;
        RECT 558.720 21.605 558.980 21.865 ;
        RECT 559.380 21.605 559.640 21.865 ;
        RECT 560.040 21.605 560.300 21.865 ;
        RECT 558.720 20.945 558.980 21.205 ;
        RECT 559.380 20.945 559.640 21.205 ;
        RECT 560.040 20.945 560.300 21.205 ;
        RECT 564.525 58.805 564.785 59.065 ;
        RECT 564.525 58.145 564.785 58.405 ;
        RECT 564.525 57.485 564.785 57.745 ;
        RECT 564.525 56.825 564.785 57.085 ;
        RECT 564.525 56.165 564.785 56.425 ;
        RECT 564.525 55.505 564.785 55.765 ;
        RECT 564.525 54.845 564.785 55.105 ;
        RECT 564.525 54.185 564.785 54.445 ;
        RECT 564.525 53.525 564.785 53.785 ;
        RECT 564.525 52.865 564.785 53.125 ;
        RECT 564.525 52.205 564.785 52.465 ;
        RECT 564.525 51.545 564.785 51.805 ;
        RECT 564.525 50.885 564.785 51.145 ;
        RECT 564.525 50.225 564.785 50.485 ;
        RECT 576.175 59.990 576.435 60.250 ;
        RECT 594.020 59.990 594.280 60.250 ;
        RECT 569.020 45.165 569.280 45.425 ;
        RECT 569.680 45.165 569.940 45.425 ;
        RECT 570.340 45.165 570.600 45.425 ;
        RECT 569.020 44.505 569.280 44.765 ;
        RECT 569.680 44.505 569.940 44.765 ;
        RECT 570.340 44.505 570.600 44.765 ;
        RECT 569.020 43.845 569.280 44.105 ;
        RECT 569.680 43.845 569.940 44.105 ;
        RECT 570.340 43.845 570.600 44.105 ;
        RECT 569.020 24.965 569.280 25.225 ;
        RECT 569.680 24.965 569.940 25.225 ;
        RECT 570.340 24.965 570.600 25.225 ;
        RECT 569.020 24.305 569.280 24.565 ;
        RECT 569.680 24.305 569.940 24.565 ;
        RECT 570.340 24.305 570.600 24.565 ;
        RECT 569.020 23.645 569.280 23.905 ;
        RECT 569.680 23.645 569.940 23.905 ;
        RECT 570.340 23.645 570.600 23.905 ;
        RECT 543.895 8.805 544.155 9.065 ;
        RECT 563.160 8.805 563.420 9.065 ;
        RECT 574.810 58.805 575.070 59.065 ;
        RECT 574.810 58.145 575.070 58.405 ;
        RECT 574.810 57.485 575.070 57.745 ;
        RECT 574.810 56.825 575.070 57.085 ;
        RECT 574.810 56.165 575.070 56.425 ;
        RECT 574.810 55.505 575.070 55.765 ;
        RECT 574.810 54.845 575.070 55.105 ;
        RECT 574.810 54.185 575.070 54.445 ;
        RECT 574.810 53.525 575.070 53.785 ;
        RECT 574.810 52.865 575.070 53.125 ;
        RECT 574.810 52.205 575.070 52.465 ;
        RECT 574.810 51.545 575.070 51.805 ;
        RECT 574.810 50.885 575.070 51.145 ;
        RECT 574.810 50.225 575.070 50.485 ;
        RECT 579.295 42.465 579.555 42.725 ;
        RECT 579.955 42.465 580.215 42.725 ;
        RECT 580.615 42.465 580.875 42.725 ;
        RECT 579.295 41.805 579.555 42.065 ;
        RECT 579.955 41.805 580.215 42.065 ;
        RECT 580.615 41.805 580.875 42.065 ;
        RECT 579.295 41.145 579.555 41.405 ;
        RECT 579.955 41.145 580.215 41.405 ;
        RECT 580.615 41.145 580.875 41.405 ;
        RECT 579.295 27.665 579.555 27.925 ;
        RECT 579.955 27.665 580.215 27.925 ;
        RECT 580.615 27.665 580.875 27.925 ;
        RECT 579.295 27.005 579.555 27.265 ;
        RECT 579.955 27.005 580.215 27.265 ;
        RECT 580.615 27.005 580.875 27.265 ;
        RECT 579.295 26.345 579.555 26.605 ;
        RECT 579.955 26.345 580.215 26.605 ;
        RECT 580.615 26.345 580.875 26.605 ;
        RECT 585.100 58.805 585.360 59.065 ;
        RECT 585.100 58.145 585.360 58.405 ;
        RECT 585.100 57.485 585.360 57.745 ;
        RECT 585.100 56.825 585.360 57.085 ;
        RECT 585.100 56.165 585.360 56.425 ;
        RECT 585.100 55.505 585.360 55.765 ;
        RECT 585.100 54.845 585.360 55.105 ;
        RECT 585.100 54.185 585.360 54.445 ;
        RECT 585.100 53.525 585.360 53.785 ;
        RECT 585.100 52.865 585.360 53.125 ;
        RECT 585.100 52.205 585.360 52.465 ;
        RECT 585.100 51.545 585.360 51.805 ;
        RECT 585.100 50.885 585.360 51.145 ;
        RECT 585.100 50.225 585.360 50.485 ;
        RECT 598.170 59.990 598.430 60.250 ;
        RECT 616.015 59.990 616.275 60.250 ;
        RECT 589.595 39.765 589.855 40.025 ;
        RECT 590.255 39.765 590.515 40.025 ;
        RECT 590.915 39.765 591.175 40.025 ;
        RECT 589.595 39.105 589.855 39.365 ;
        RECT 590.255 39.105 590.515 39.365 ;
        RECT 590.915 39.105 591.175 39.365 ;
        RECT 589.595 38.445 589.855 38.705 ;
        RECT 590.255 38.445 590.515 38.705 ;
        RECT 590.915 38.445 591.175 38.705 ;
        RECT 589.595 30.365 589.855 30.625 ;
        RECT 590.255 30.365 590.515 30.625 ;
        RECT 590.915 30.365 591.175 30.625 ;
        RECT 589.595 29.705 589.855 29.965 ;
        RECT 590.255 29.705 590.515 29.965 ;
        RECT 590.915 29.705 591.175 29.965 ;
        RECT 589.595 29.045 589.855 29.305 ;
        RECT 590.255 29.045 590.515 29.305 ;
        RECT 590.915 29.045 591.175 29.305 ;
        RECT 565.890 8.805 566.150 9.065 ;
        RECT 583.735 8.805 583.995 9.065 ;
        RECT 595.385 58.805 595.645 59.065 ;
        RECT 595.385 58.145 595.645 58.405 ;
        RECT 595.385 57.485 595.645 57.745 ;
        RECT 595.385 56.825 595.645 57.085 ;
        RECT 595.385 56.165 595.645 56.425 ;
        RECT 595.385 55.505 595.645 55.765 ;
        RECT 595.385 54.845 595.645 55.105 ;
        RECT 595.385 54.185 595.645 54.445 ;
        RECT 595.385 53.525 595.645 53.785 ;
        RECT 595.385 52.865 595.645 53.125 ;
        RECT 595.385 52.205 595.645 52.465 ;
        RECT 595.385 51.545 595.645 51.805 ;
        RECT 595.385 50.885 595.645 51.145 ;
        RECT 595.385 50.225 595.645 50.485 ;
        RECT 596.805 58.805 597.065 59.065 ;
        RECT 596.805 58.145 597.065 58.405 ;
        RECT 596.805 57.485 597.065 57.745 ;
        RECT 596.805 56.825 597.065 57.085 ;
        RECT 596.805 56.165 597.065 56.425 ;
        RECT 596.805 55.505 597.065 55.765 ;
        RECT 596.805 54.845 597.065 55.105 ;
        RECT 596.805 54.185 597.065 54.445 ;
        RECT 596.805 53.525 597.065 53.785 ;
        RECT 596.805 52.865 597.065 53.125 ;
        RECT 596.805 52.205 597.065 52.465 ;
        RECT 596.805 51.545 597.065 51.805 ;
        RECT 596.805 50.885 597.065 51.145 ;
        RECT 596.805 50.225 597.065 50.485 ;
        RECT 601.290 47.865 601.550 48.125 ;
        RECT 601.950 47.865 602.210 48.125 ;
        RECT 602.610 47.865 602.870 48.125 ;
        RECT 601.290 47.205 601.550 47.465 ;
        RECT 601.950 47.205 602.210 47.465 ;
        RECT 602.610 47.205 602.870 47.465 ;
        RECT 601.290 46.545 601.550 46.805 ;
        RECT 601.950 46.545 602.210 46.805 ;
        RECT 602.610 46.545 602.870 46.805 ;
        RECT 601.290 22.265 601.550 22.525 ;
        RECT 601.950 22.265 602.210 22.525 ;
        RECT 602.610 22.265 602.870 22.525 ;
        RECT 601.290 21.605 601.550 21.865 ;
        RECT 601.950 21.605 602.210 21.865 ;
        RECT 602.610 21.605 602.870 21.865 ;
        RECT 601.290 20.945 601.550 21.205 ;
        RECT 601.950 20.945 602.210 21.205 ;
        RECT 602.610 20.945 602.870 21.205 ;
        RECT 607.095 58.805 607.355 59.065 ;
        RECT 607.095 58.145 607.355 58.405 ;
        RECT 607.095 57.485 607.355 57.745 ;
        RECT 607.095 56.825 607.355 57.085 ;
        RECT 607.095 56.165 607.355 56.425 ;
        RECT 607.095 55.505 607.355 55.765 ;
        RECT 607.095 54.845 607.355 55.105 ;
        RECT 607.095 54.185 607.355 54.445 ;
        RECT 607.095 53.525 607.355 53.785 ;
        RECT 607.095 52.865 607.355 53.125 ;
        RECT 607.095 52.205 607.355 52.465 ;
        RECT 607.095 51.545 607.355 51.805 ;
        RECT 607.095 50.885 607.355 51.145 ;
        RECT 607.095 50.225 607.355 50.485 ;
        RECT 618.745 59.990 619.005 60.250 ;
        RECT 636.590 59.990 636.850 60.250 ;
        RECT 611.590 45.165 611.850 45.425 ;
        RECT 612.250 45.165 612.510 45.425 ;
        RECT 612.910 45.165 613.170 45.425 ;
        RECT 611.590 44.505 611.850 44.765 ;
        RECT 612.250 44.505 612.510 44.765 ;
        RECT 612.910 44.505 613.170 44.765 ;
        RECT 611.590 43.845 611.850 44.105 ;
        RECT 612.250 43.845 612.510 44.105 ;
        RECT 612.910 43.845 613.170 44.105 ;
        RECT 611.590 24.965 611.850 25.225 ;
        RECT 612.250 24.965 612.510 25.225 ;
        RECT 612.910 24.965 613.170 25.225 ;
        RECT 611.590 24.305 611.850 24.565 ;
        RECT 612.250 24.305 612.510 24.565 ;
        RECT 612.910 24.305 613.170 24.565 ;
        RECT 611.590 23.645 611.850 23.905 ;
        RECT 612.250 23.645 612.510 23.905 ;
        RECT 612.910 23.645 613.170 23.905 ;
        RECT 586.465 8.805 586.725 9.065 ;
        RECT 605.730 8.805 605.990 9.065 ;
        RECT 617.380 58.805 617.640 59.065 ;
        RECT 617.380 58.145 617.640 58.405 ;
        RECT 617.380 57.485 617.640 57.745 ;
        RECT 617.380 56.825 617.640 57.085 ;
        RECT 617.380 56.165 617.640 56.425 ;
        RECT 617.380 55.505 617.640 55.765 ;
        RECT 617.380 54.845 617.640 55.105 ;
        RECT 617.380 54.185 617.640 54.445 ;
        RECT 617.380 53.525 617.640 53.785 ;
        RECT 617.380 52.865 617.640 53.125 ;
        RECT 617.380 52.205 617.640 52.465 ;
        RECT 617.380 51.545 617.640 51.805 ;
        RECT 617.380 50.885 617.640 51.145 ;
        RECT 617.380 50.225 617.640 50.485 ;
        RECT 621.865 42.465 622.125 42.725 ;
        RECT 622.525 42.465 622.785 42.725 ;
        RECT 623.185 42.465 623.445 42.725 ;
        RECT 621.865 41.805 622.125 42.065 ;
        RECT 622.525 41.805 622.785 42.065 ;
        RECT 623.185 41.805 623.445 42.065 ;
        RECT 621.865 41.145 622.125 41.405 ;
        RECT 622.525 41.145 622.785 41.405 ;
        RECT 623.185 41.145 623.445 41.405 ;
        RECT 621.865 27.665 622.125 27.925 ;
        RECT 622.525 27.665 622.785 27.925 ;
        RECT 623.185 27.665 623.445 27.925 ;
        RECT 621.865 27.005 622.125 27.265 ;
        RECT 622.525 27.005 622.785 27.265 ;
        RECT 623.185 27.005 623.445 27.265 ;
        RECT 621.865 26.345 622.125 26.605 ;
        RECT 622.525 26.345 622.785 26.605 ;
        RECT 623.185 26.345 623.445 26.605 ;
        RECT 627.670 58.805 627.930 59.065 ;
        RECT 627.670 58.145 627.930 58.405 ;
        RECT 627.670 57.485 627.930 57.745 ;
        RECT 627.670 56.825 627.930 57.085 ;
        RECT 627.670 56.165 627.930 56.425 ;
        RECT 627.670 55.505 627.930 55.765 ;
        RECT 627.670 54.845 627.930 55.105 ;
        RECT 627.670 54.185 627.930 54.445 ;
        RECT 627.670 53.525 627.930 53.785 ;
        RECT 627.670 52.865 627.930 53.125 ;
        RECT 627.670 52.205 627.930 52.465 ;
        RECT 627.670 51.545 627.930 51.805 ;
        RECT 627.670 50.885 627.930 51.145 ;
        RECT 627.670 50.225 627.930 50.485 ;
        RECT 640.740 59.990 641.000 60.250 ;
        RECT 658.585 59.990 658.845 60.250 ;
        RECT 632.165 39.765 632.425 40.025 ;
        RECT 632.825 39.765 633.085 40.025 ;
        RECT 633.485 39.765 633.745 40.025 ;
        RECT 632.165 39.105 632.425 39.365 ;
        RECT 632.825 39.105 633.085 39.365 ;
        RECT 633.485 39.105 633.745 39.365 ;
        RECT 632.165 38.445 632.425 38.705 ;
        RECT 632.825 38.445 633.085 38.705 ;
        RECT 633.485 38.445 633.745 38.705 ;
        RECT 632.165 30.365 632.425 30.625 ;
        RECT 632.825 30.365 633.085 30.625 ;
        RECT 633.485 30.365 633.745 30.625 ;
        RECT 632.165 29.705 632.425 29.965 ;
        RECT 632.825 29.705 633.085 29.965 ;
        RECT 633.485 29.705 633.745 29.965 ;
        RECT 632.165 29.045 632.425 29.305 ;
        RECT 632.825 29.045 633.085 29.305 ;
        RECT 633.485 29.045 633.745 29.305 ;
        RECT 608.460 8.805 608.720 9.065 ;
        RECT 626.305 8.805 626.565 9.065 ;
        RECT 637.955 58.805 638.215 59.065 ;
        RECT 637.955 58.145 638.215 58.405 ;
        RECT 637.955 57.485 638.215 57.745 ;
        RECT 637.955 56.825 638.215 57.085 ;
        RECT 637.955 56.165 638.215 56.425 ;
        RECT 637.955 55.505 638.215 55.765 ;
        RECT 637.955 54.845 638.215 55.105 ;
        RECT 637.955 54.185 638.215 54.445 ;
        RECT 637.955 53.525 638.215 53.785 ;
        RECT 637.955 52.865 638.215 53.125 ;
        RECT 637.955 52.205 638.215 52.465 ;
        RECT 637.955 51.545 638.215 51.805 ;
        RECT 637.955 50.885 638.215 51.145 ;
        RECT 637.955 50.225 638.215 50.485 ;
        RECT 639.375 58.805 639.635 59.065 ;
        RECT 639.375 58.145 639.635 58.405 ;
        RECT 639.375 57.485 639.635 57.745 ;
        RECT 639.375 56.825 639.635 57.085 ;
        RECT 639.375 56.165 639.635 56.425 ;
        RECT 639.375 55.505 639.635 55.765 ;
        RECT 639.375 54.845 639.635 55.105 ;
        RECT 639.375 54.185 639.635 54.445 ;
        RECT 639.375 53.525 639.635 53.785 ;
        RECT 639.375 52.865 639.635 53.125 ;
        RECT 639.375 52.205 639.635 52.465 ;
        RECT 639.375 51.545 639.635 51.805 ;
        RECT 639.375 50.885 639.635 51.145 ;
        RECT 639.375 50.225 639.635 50.485 ;
        RECT 643.860 47.865 644.120 48.125 ;
        RECT 644.520 47.865 644.780 48.125 ;
        RECT 645.180 47.865 645.440 48.125 ;
        RECT 643.860 47.205 644.120 47.465 ;
        RECT 644.520 47.205 644.780 47.465 ;
        RECT 645.180 47.205 645.440 47.465 ;
        RECT 643.860 46.545 644.120 46.805 ;
        RECT 644.520 46.545 644.780 46.805 ;
        RECT 645.180 46.545 645.440 46.805 ;
        RECT 643.860 22.265 644.120 22.525 ;
        RECT 644.520 22.265 644.780 22.525 ;
        RECT 645.180 22.265 645.440 22.525 ;
        RECT 643.860 21.605 644.120 21.865 ;
        RECT 644.520 21.605 644.780 21.865 ;
        RECT 645.180 21.605 645.440 21.865 ;
        RECT 643.860 20.945 644.120 21.205 ;
        RECT 644.520 20.945 644.780 21.205 ;
        RECT 645.180 20.945 645.440 21.205 ;
        RECT 649.665 58.805 649.925 59.065 ;
        RECT 649.665 58.145 649.925 58.405 ;
        RECT 649.665 57.485 649.925 57.745 ;
        RECT 649.665 56.825 649.925 57.085 ;
        RECT 649.665 56.165 649.925 56.425 ;
        RECT 649.665 55.505 649.925 55.765 ;
        RECT 649.665 54.845 649.925 55.105 ;
        RECT 649.665 54.185 649.925 54.445 ;
        RECT 649.665 53.525 649.925 53.785 ;
        RECT 649.665 52.865 649.925 53.125 ;
        RECT 649.665 52.205 649.925 52.465 ;
        RECT 649.665 51.545 649.925 51.805 ;
        RECT 649.665 50.885 649.925 51.145 ;
        RECT 649.665 50.225 649.925 50.485 ;
        RECT 661.315 59.990 661.575 60.250 ;
        RECT 679.160 59.990 679.420 60.250 ;
        RECT 654.160 45.165 654.420 45.425 ;
        RECT 654.820 45.165 655.080 45.425 ;
        RECT 655.480 45.165 655.740 45.425 ;
        RECT 654.160 44.505 654.420 44.765 ;
        RECT 654.820 44.505 655.080 44.765 ;
        RECT 655.480 44.505 655.740 44.765 ;
        RECT 654.160 43.845 654.420 44.105 ;
        RECT 654.820 43.845 655.080 44.105 ;
        RECT 655.480 43.845 655.740 44.105 ;
        RECT 654.160 24.965 654.420 25.225 ;
        RECT 654.820 24.965 655.080 25.225 ;
        RECT 655.480 24.965 655.740 25.225 ;
        RECT 654.160 24.305 654.420 24.565 ;
        RECT 654.820 24.305 655.080 24.565 ;
        RECT 655.480 24.305 655.740 24.565 ;
        RECT 654.160 23.645 654.420 23.905 ;
        RECT 654.820 23.645 655.080 23.905 ;
        RECT 655.480 23.645 655.740 23.905 ;
        RECT 629.035 8.805 629.295 9.065 ;
        RECT 648.300 8.805 648.560 9.065 ;
        RECT 659.950 58.805 660.210 59.065 ;
        RECT 659.950 58.145 660.210 58.405 ;
        RECT 659.950 57.485 660.210 57.745 ;
        RECT 659.950 56.825 660.210 57.085 ;
        RECT 659.950 56.165 660.210 56.425 ;
        RECT 659.950 55.505 660.210 55.765 ;
        RECT 659.950 54.845 660.210 55.105 ;
        RECT 659.950 54.185 660.210 54.445 ;
        RECT 659.950 53.525 660.210 53.785 ;
        RECT 659.950 52.865 660.210 53.125 ;
        RECT 659.950 52.205 660.210 52.465 ;
        RECT 659.950 51.545 660.210 51.805 ;
        RECT 659.950 50.885 660.210 51.145 ;
        RECT 659.950 50.225 660.210 50.485 ;
        RECT 664.435 42.465 664.695 42.725 ;
        RECT 665.095 42.465 665.355 42.725 ;
        RECT 665.755 42.465 666.015 42.725 ;
        RECT 664.435 41.805 664.695 42.065 ;
        RECT 665.095 41.805 665.355 42.065 ;
        RECT 665.755 41.805 666.015 42.065 ;
        RECT 664.435 41.145 664.695 41.405 ;
        RECT 665.095 41.145 665.355 41.405 ;
        RECT 665.755 41.145 666.015 41.405 ;
        RECT 664.435 27.665 664.695 27.925 ;
        RECT 665.095 27.665 665.355 27.925 ;
        RECT 665.755 27.665 666.015 27.925 ;
        RECT 664.435 27.005 664.695 27.265 ;
        RECT 665.095 27.005 665.355 27.265 ;
        RECT 665.755 27.005 666.015 27.265 ;
        RECT 664.435 26.345 664.695 26.605 ;
        RECT 665.095 26.345 665.355 26.605 ;
        RECT 665.755 26.345 666.015 26.605 ;
        RECT 670.240 58.805 670.500 59.065 ;
        RECT 670.240 58.145 670.500 58.405 ;
        RECT 670.240 57.485 670.500 57.745 ;
        RECT 670.240 56.825 670.500 57.085 ;
        RECT 670.240 56.165 670.500 56.425 ;
        RECT 670.240 55.505 670.500 55.765 ;
        RECT 670.240 54.845 670.500 55.105 ;
        RECT 670.240 54.185 670.500 54.445 ;
        RECT 670.240 53.525 670.500 53.785 ;
        RECT 670.240 52.865 670.500 53.125 ;
        RECT 670.240 52.205 670.500 52.465 ;
        RECT 670.240 51.545 670.500 51.805 ;
        RECT 670.240 50.885 670.500 51.145 ;
        RECT 670.240 50.225 670.500 50.485 ;
        RECT 674.735 39.765 674.995 40.025 ;
        RECT 675.395 39.765 675.655 40.025 ;
        RECT 676.055 39.765 676.315 40.025 ;
        RECT 674.735 39.105 674.995 39.365 ;
        RECT 675.395 39.105 675.655 39.365 ;
        RECT 676.055 39.105 676.315 39.365 ;
        RECT 674.735 38.445 674.995 38.705 ;
        RECT 675.395 38.445 675.655 38.705 ;
        RECT 676.055 38.445 676.315 38.705 ;
        RECT 674.735 30.365 674.995 30.625 ;
        RECT 675.395 30.365 675.655 30.625 ;
        RECT 676.055 30.365 676.315 30.625 ;
        RECT 674.735 29.705 674.995 29.965 ;
        RECT 675.395 29.705 675.655 29.965 ;
        RECT 676.055 29.705 676.315 29.965 ;
        RECT 674.735 29.045 674.995 29.305 ;
        RECT 675.395 29.045 675.655 29.305 ;
        RECT 676.055 29.045 676.315 29.305 ;
        RECT 651.030 8.805 651.290 9.065 ;
        RECT 668.875 8.805 669.135 9.065 ;
        RECT 680.525 58.805 680.785 59.065 ;
        RECT 680.525 58.145 680.785 58.405 ;
        RECT 680.525 57.485 680.785 57.745 ;
        RECT 680.525 56.825 680.785 57.085 ;
        RECT 680.525 56.165 680.785 56.425 ;
        RECT 680.525 55.505 680.785 55.765 ;
        RECT 680.525 54.845 680.785 55.105 ;
        RECT 680.525 54.185 680.785 54.445 ;
        RECT 680.525 53.525 680.785 53.785 ;
        RECT 680.525 52.865 680.785 53.125 ;
        RECT 680.525 52.205 680.785 52.465 ;
        RECT 680.525 51.545 680.785 51.805 ;
        RECT 680.525 50.885 680.785 51.145 ;
        RECT 680.525 50.225 680.785 50.485 ;
        RECT 682.370 55.175 682.630 55.435 ;
        RECT 682.370 54.515 682.630 54.775 ;
        RECT 682.370 53.855 682.630 54.115 ;
        RECT 682.370 53.195 682.630 53.455 ;
        RECT 682.370 52.535 682.630 52.795 ;
        RECT 682.370 51.875 682.630 52.135 ;
        RECT 682.370 51.215 682.630 51.475 ;
        RECT 682.370 50.555 682.630 50.815 ;
        RECT 682.370 18.175 682.630 18.435 ;
        RECT 682.370 17.515 682.630 17.775 ;
        RECT 682.370 16.855 682.630 17.115 ;
        RECT 682.370 16.195 682.630 16.455 ;
        RECT 682.370 15.535 682.630 15.795 ;
        RECT 682.370 14.875 682.630 15.135 ;
        RECT 682.370 14.215 682.630 14.475 ;
        RECT 682.370 13.555 682.630 13.815 ;
        RECT 682.370 12.895 682.630 13.155 ;
        RECT 682.370 12.235 682.630 12.495 ;
        RECT 682.370 11.575 682.630 11.835 ;
        RECT 682.370 10.915 682.630 11.175 ;
        RECT 682.370 10.255 682.630 10.515 ;
        RECT 682.370 9.595 682.630 9.855 ;
        RECT 671.605 8.805 671.865 9.065 ;
        RECT 682.370 8.935 682.630 9.195 ;
        RECT 684.155 55.175 684.415 55.435 ;
        RECT 687.010 55.175 687.270 55.435 ;
        RECT 684.155 54.515 684.415 54.775 ;
        RECT 687.010 54.515 687.270 54.775 ;
        RECT 684.155 53.855 684.415 54.115 ;
        RECT 687.010 53.855 687.270 54.115 ;
        RECT 684.155 53.195 684.415 53.455 ;
        RECT 687.010 53.195 687.270 53.455 ;
        RECT 684.155 52.535 684.415 52.795 ;
        RECT 687.010 52.535 687.270 52.795 ;
        RECT 684.155 51.875 684.415 52.135 ;
        RECT 687.010 51.875 687.270 52.135 ;
        RECT 684.155 51.215 684.415 51.475 ;
        RECT 687.010 51.215 687.270 51.475 ;
        RECT 684.155 50.555 684.415 50.815 ;
        RECT 687.010 50.555 687.270 50.815 ;
        RECT 683.130 47.865 683.390 48.125 ;
        RECT 683.130 47.205 683.390 47.465 ;
        RECT 683.130 46.545 683.390 46.805 ;
        RECT 684.155 18.175 684.415 18.435 ;
        RECT 687.010 18.175 687.270 18.435 ;
        RECT 684.155 17.515 684.415 17.775 ;
        RECT 687.010 17.515 687.270 17.775 ;
        RECT 684.155 16.855 684.415 17.115 ;
        RECT 687.010 16.855 687.270 17.115 ;
        RECT 684.155 16.195 684.415 16.455 ;
        RECT 687.010 16.195 687.270 16.455 ;
        RECT 684.155 15.535 684.415 15.795 ;
        RECT 687.010 15.535 687.270 15.795 ;
        RECT 684.155 14.875 684.415 15.135 ;
        RECT 687.010 14.875 687.270 15.135 ;
        RECT 684.155 14.215 684.415 14.475 ;
        RECT 687.010 14.215 687.270 14.475 ;
        RECT 684.155 13.555 684.415 13.815 ;
        RECT 687.010 13.555 687.270 13.815 ;
        RECT 684.155 12.895 684.415 13.155 ;
        RECT 687.010 12.895 687.270 13.155 ;
        RECT 684.155 12.235 684.415 12.495 ;
        RECT 687.010 12.235 687.270 12.495 ;
        RECT 684.155 11.575 684.415 11.835 ;
        RECT 687.010 11.575 687.270 11.835 ;
        RECT 684.155 10.915 684.415 11.175 ;
        RECT 687.010 10.915 687.270 11.175 ;
        RECT 684.155 10.255 684.415 10.515 ;
        RECT 687.010 10.255 687.270 10.515 ;
        RECT 684.155 9.595 684.415 9.855 ;
        RECT 687.010 9.595 687.270 9.855 ;
        RECT 684.155 8.935 684.415 9.195 ;
        RECT 687.010 8.935 687.270 9.195 ;
        RECT 688.795 55.175 689.055 55.435 ;
        RECT 691.650 55.175 691.910 55.435 ;
        RECT 688.795 54.515 689.055 54.775 ;
        RECT 691.650 54.515 691.910 54.775 ;
        RECT 688.795 53.855 689.055 54.115 ;
        RECT 691.650 53.855 691.910 54.115 ;
        RECT 688.795 53.195 689.055 53.455 ;
        RECT 691.650 53.195 691.910 53.455 ;
        RECT 688.795 52.535 689.055 52.795 ;
        RECT 691.650 52.535 691.910 52.795 ;
        RECT 688.795 51.875 689.055 52.135 ;
        RECT 691.650 51.875 691.910 52.135 ;
        RECT 688.795 51.215 689.055 51.475 ;
        RECT 691.650 51.215 691.910 51.475 ;
        RECT 688.795 50.555 689.055 50.815 ;
        RECT 691.650 50.555 691.910 50.815 ;
        RECT 687.770 22.265 688.030 22.525 ;
        RECT 687.770 21.605 688.030 21.865 ;
        RECT 687.770 20.945 688.030 21.205 ;
        RECT 688.795 18.175 689.055 18.435 ;
        RECT 691.650 18.175 691.910 18.435 ;
        RECT 688.795 17.515 689.055 17.775 ;
        RECT 691.650 17.515 691.910 17.775 ;
        RECT 688.795 16.855 689.055 17.115 ;
        RECT 691.650 16.855 691.910 17.115 ;
        RECT 688.795 16.195 689.055 16.455 ;
        RECT 691.650 16.195 691.910 16.455 ;
        RECT 688.795 15.535 689.055 15.795 ;
        RECT 691.650 15.535 691.910 15.795 ;
        RECT 688.795 14.875 689.055 15.135 ;
        RECT 691.650 14.875 691.910 15.135 ;
        RECT 688.795 14.215 689.055 14.475 ;
        RECT 691.650 14.215 691.910 14.475 ;
        RECT 688.795 13.555 689.055 13.815 ;
        RECT 691.650 13.555 691.910 13.815 ;
        RECT 688.795 12.895 689.055 13.155 ;
        RECT 691.650 12.895 691.910 13.155 ;
        RECT 688.795 12.235 689.055 12.495 ;
        RECT 691.650 12.235 691.910 12.495 ;
        RECT 688.795 11.575 689.055 11.835 ;
        RECT 691.650 11.575 691.910 11.835 ;
        RECT 688.795 10.915 689.055 11.175 ;
        RECT 691.650 10.915 691.910 11.175 ;
        RECT 688.795 10.255 689.055 10.515 ;
        RECT 691.650 10.255 691.910 10.515 ;
        RECT 688.795 9.595 689.055 9.855 ;
        RECT 691.650 9.595 691.910 9.855 ;
        RECT 688.795 8.935 689.055 9.195 ;
        RECT 691.650 8.935 691.910 9.195 ;
        RECT 693.435 55.175 693.695 55.435 ;
        RECT 696.290 55.175 696.550 55.435 ;
        RECT 693.435 54.515 693.695 54.775 ;
        RECT 696.290 54.515 696.550 54.775 ;
        RECT 693.435 53.855 693.695 54.115 ;
        RECT 696.290 53.855 696.550 54.115 ;
        RECT 693.435 53.195 693.695 53.455 ;
        RECT 696.290 53.195 696.550 53.455 ;
        RECT 693.435 52.535 693.695 52.795 ;
        RECT 696.290 52.535 696.550 52.795 ;
        RECT 693.435 51.875 693.695 52.135 ;
        RECT 696.290 51.875 696.550 52.135 ;
        RECT 693.435 51.215 693.695 51.475 ;
        RECT 696.290 51.215 696.550 51.475 ;
        RECT 693.435 50.555 693.695 50.815 ;
        RECT 696.290 50.555 696.550 50.815 ;
        RECT 692.410 24.965 692.670 25.225 ;
        RECT 692.410 24.305 692.670 24.565 ;
        RECT 692.410 23.645 692.670 23.905 ;
        RECT 693.435 18.175 693.695 18.435 ;
        RECT 696.290 18.175 696.550 18.435 ;
        RECT 693.435 17.515 693.695 17.775 ;
        RECT 696.290 17.515 696.550 17.775 ;
        RECT 693.435 16.855 693.695 17.115 ;
        RECT 696.290 16.855 696.550 17.115 ;
        RECT 693.435 16.195 693.695 16.455 ;
        RECT 696.290 16.195 696.550 16.455 ;
        RECT 693.435 15.535 693.695 15.795 ;
        RECT 696.290 15.535 696.550 15.795 ;
        RECT 693.435 14.875 693.695 15.135 ;
        RECT 696.290 14.875 696.550 15.135 ;
        RECT 693.435 14.215 693.695 14.475 ;
        RECT 696.290 14.215 696.550 14.475 ;
        RECT 693.435 13.555 693.695 13.815 ;
        RECT 696.290 13.555 696.550 13.815 ;
        RECT 693.435 12.895 693.695 13.155 ;
        RECT 696.290 12.895 696.550 13.155 ;
        RECT 693.435 12.235 693.695 12.495 ;
        RECT 696.290 12.235 696.550 12.495 ;
        RECT 693.435 11.575 693.695 11.835 ;
        RECT 696.290 11.575 696.550 11.835 ;
        RECT 693.435 10.915 693.695 11.175 ;
        RECT 696.290 10.915 696.550 11.175 ;
        RECT 693.435 10.255 693.695 10.515 ;
        RECT 696.290 10.255 696.550 10.515 ;
        RECT 693.435 9.595 693.695 9.855 ;
        RECT 696.290 9.595 696.550 9.855 ;
        RECT 693.435 8.935 693.695 9.195 ;
        RECT 696.290 8.935 696.550 9.195 ;
        RECT 698.075 55.175 698.335 55.435 ;
        RECT 700.930 55.175 701.190 55.435 ;
        RECT 698.075 54.515 698.335 54.775 ;
        RECT 700.930 54.515 701.190 54.775 ;
        RECT 698.075 53.855 698.335 54.115 ;
        RECT 700.930 53.855 701.190 54.115 ;
        RECT 698.075 53.195 698.335 53.455 ;
        RECT 700.930 53.195 701.190 53.455 ;
        RECT 698.075 52.535 698.335 52.795 ;
        RECT 700.930 52.535 701.190 52.795 ;
        RECT 698.075 51.875 698.335 52.135 ;
        RECT 700.930 51.875 701.190 52.135 ;
        RECT 698.075 51.215 698.335 51.475 ;
        RECT 700.930 51.215 701.190 51.475 ;
        RECT 698.075 50.555 698.335 50.815 ;
        RECT 700.930 50.555 701.190 50.815 ;
        RECT 697.050 45.165 697.310 45.425 ;
        RECT 697.050 44.505 697.310 44.765 ;
        RECT 697.050 43.845 697.310 44.105 ;
        RECT 698.075 18.175 698.335 18.435 ;
        RECT 700.930 18.175 701.190 18.435 ;
        RECT 698.075 17.515 698.335 17.775 ;
        RECT 700.930 17.515 701.190 17.775 ;
        RECT 698.075 16.855 698.335 17.115 ;
        RECT 700.930 16.855 701.190 17.115 ;
        RECT 698.075 16.195 698.335 16.455 ;
        RECT 700.930 16.195 701.190 16.455 ;
        RECT 698.075 15.535 698.335 15.795 ;
        RECT 700.930 15.535 701.190 15.795 ;
        RECT 698.075 14.875 698.335 15.135 ;
        RECT 700.930 14.875 701.190 15.135 ;
        RECT 698.075 14.215 698.335 14.475 ;
        RECT 700.930 14.215 701.190 14.475 ;
        RECT 698.075 13.555 698.335 13.815 ;
        RECT 700.930 13.555 701.190 13.815 ;
        RECT 698.075 12.895 698.335 13.155 ;
        RECT 700.930 12.895 701.190 13.155 ;
        RECT 698.075 12.235 698.335 12.495 ;
        RECT 700.930 12.235 701.190 12.495 ;
        RECT 698.075 11.575 698.335 11.835 ;
        RECT 700.930 11.575 701.190 11.835 ;
        RECT 698.075 10.915 698.335 11.175 ;
        RECT 700.930 10.915 701.190 11.175 ;
        RECT 698.075 10.255 698.335 10.515 ;
        RECT 700.930 10.255 701.190 10.515 ;
        RECT 698.075 9.595 698.335 9.855 ;
        RECT 700.930 9.595 701.190 9.855 ;
        RECT 698.075 8.935 698.335 9.195 ;
        RECT 700.930 8.935 701.190 9.195 ;
        RECT 702.715 55.175 702.975 55.435 ;
        RECT 705.570 55.175 705.830 55.435 ;
        RECT 702.715 54.515 702.975 54.775 ;
        RECT 705.570 54.515 705.830 54.775 ;
        RECT 702.715 53.855 702.975 54.115 ;
        RECT 705.570 53.855 705.830 54.115 ;
        RECT 702.715 53.195 702.975 53.455 ;
        RECT 705.570 53.195 705.830 53.455 ;
        RECT 702.715 52.535 702.975 52.795 ;
        RECT 705.570 52.535 705.830 52.795 ;
        RECT 702.715 51.875 702.975 52.135 ;
        RECT 705.570 51.875 705.830 52.135 ;
        RECT 702.715 51.215 702.975 51.475 ;
        RECT 705.570 51.215 705.830 51.475 ;
        RECT 702.715 50.555 702.975 50.815 ;
        RECT 705.570 50.555 705.830 50.815 ;
        RECT 701.690 42.465 701.950 42.725 ;
        RECT 701.690 41.805 701.950 42.065 ;
        RECT 701.690 41.145 701.950 41.405 ;
        RECT 702.715 18.175 702.975 18.435 ;
        RECT 705.570 18.175 705.830 18.435 ;
        RECT 702.715 17.515 702.975 17.775 ;
        RECT 705.570 17.515 705.830 17.775 ;
        RECT 702.715 16.855 702.975 17.115 ;
        RECT 705.570 16.855 705.830 17.115 ;
        RECT 702.715 16.195 702.975 16.455 ;
        RECT 705.570 16.195 705.830 16.455 ;
        RECT 702.715 15.535 702.975 15.795 ;
        RECT 705.570 15.535 705.830 15.795 ;
        RECT 702.715 14.875 702.975 15.135 ;
        RECT 705.570 14.875 705.830 15.135 ;
        RECT 702.715 14.215 702.975 14.475 ;
        RECT 705.570 14.215 705.830 14.475 ;
        RECT 702.715 13.555 702.975 13.815 ;
        RECT 705.570 13.555 705.830 13.815 ;
        RECT 702.715 12.895 702.975 13.155 ;
        RECT 705.570 12.895 705.830 13.155 ;
        RECT 702.715 12.235 702.975 12.495 ;
        RECT 705.570 12.235 705.830 12.495 ;
        RECT 702.715 11.575 702.975 11.835 ;
        RECT 705.570 11.575 705.830 11.835 ;
        RECT 702.715 10.915 702.975 11.175 ;
        RECT 705.570 10.915 705.830 11.175 ;
        RECT 702.715 10.255 702.975 10.515 ;
        RECT 705.570 10.255 705.830 10.515 ;
        RECT 702.715 9.595 702.975 9.855 ;
        RECT 705.570 9.595 705.830 9.855 ;
        RECT 702.715 8.935 702.975 9.195 ;
        RECT 705.570 8.935 705.830 9.195 ;
        RECT 707.355 55.175 707.615 55.435 ;
        RECT 710.210 55.175 710.470 55.435 ;
        RECT 707.355 54.515 707.615 54.775 ;
        RECT 710.210 54.515 710.470 54.775 ;
        RECT 707.355 53.855 707.615 54.115 ;
        RECT 710.210 53.855 710.470 54.115 ;
        RECT 707.355 53.195 707.615 53.455 ;
        RECT 710.210 53.195 710.470 53.455 ;
        RECT 707.355 52.535 707.615 52.795 ;
        RECT 710.210 52.535 710.470 52.795 ;
        RECT 707.355 51.875 707.615 52.135 ;
        RECT 710.210 51.875 710.470 52.135 ;
        RECT 707.355 51.215 707.615 51.475 ;
        RECT 710.210 51.215 710.470 51.475 ;
        RECT 707.355 50.555 707.615 50.815 ;
        RECT 710.210 50.555 710.470 50.815 ;
        RECT 706.330 27.665 706.590 27.925 ;
        RECT 706.330 27.005 706.590 27.265 ;
        RECT 706.330 26.345 706.590 26.605 ;
        RECT 707.355 18.175 707.615 18.435 ;
        RECT 710.210 18.175 710.470 18.435 ;
        RECT 707.355 17.515 707.615 17.775 ;
        RECT 710.210 17.515 710.470 17.775 ;
        RECT 707.355 16.855 707.615 17.115 ;
        RECT 710.210 16.855 710.470 17.115 ;
        RECT 707.355 16.195 707.615 16.455 ;
        RECT 710.210 16.195 710.470 16.455 ;
        RECT 707.355 15.535 707.615 15.795 ;
        RECT 710.210 15.535 710.470 15.795 ;
        RECT 707.355 14.875 707.615 15.135 ;
        RECT 710.210 14.875 710.470 15.135 ;
        RECT 707.355 14.215 707.615 14.475 ;
        RECT 710.210 14.215 710.470 14.475 ;
        RECT 707.355 13.555 707.615 13.815 ;
        RECT 710.210 13.555 710.470 13.815 ;
        RECT 707.355 12.895 707.615 13.155 ;
        RECT 710.210 12.895 710.470 13.155 ;
        RECT 707.355 12.235 707.615 12.495 ;
        RECT 710.210 12.235 710.470 12.495 ;
        RECT 707.355 11.575 707.615 11.835 ;
        RECT 710.210 11.575 710.470 11.835 ;
        RECT 707.355 10.915 707.615 11.175 ;
        RECT 710.210 10.915 710.470 11.175 ;
        RECT 707.355 10.255 707.615 10.515 ;
        RECT 710.210 10.255 710.470 10.515 ;
        RECT 707.355 9.595 707.615 9.855 ;
        RECT 710.210 9.595 710.470 9.855 ;
        RECT 707.355 8.935 707.615 9.195 ;
        RECT 710.210 8.935 710.470 9.195 ;
        RECT 711.995 55.175 712.255 55.435 ;
        RECT 714.850 55.175 715.110 55.435 ;
        RECT 711.995 54.515 712.255 54.775 ;
        RECT 714.850 54.515 715.110 54.775 ;
        RECT 711.995 53.855 712.255 54.115 ;
        RECT 714.850 53.855 715.110 54.115 ;
        RECT 711.995 53.195 712.255 53.455 ;
        RECT 714.850 53.195 715.110 53.455 ;
        RECT 711.995 52.535 712.255 52.795 ;
        RECT 714.850 52.535 715.110 52.795 ;
        RECT 711.995 51.875 712.255 52.135 ;
        RECT 714.850 51.875 715.110 52.135 ;
        RECT 711.995 51.215 712.255 51.475 ;
        RECT 714.850 51.215 715.110 51.475 ;
        RECT 711.995 50.555 712.255 50.815 ;
        RECT 714.850 50.555 715.110 50.815 ;
        RECT 710.970 30.365 711.230 30.625 ;
        RECT 710.970 29.705 711.230 29.965 ;
        RECT 710.970 29.045 711.230 29.305 ;
        RECT 711.995 18.175 712.255 18.435 ;
        RECT 714.850 18.175 715.110 18.435 ;
        RECT 711.995 17.515 712.255 17.775 ;
        RECT 714.850 17.515 715.110 17.775 ;
        RECT 711.995 16.855 712.255 17.115 ;
        RECT 714.850 16.855 715.110 17.115 ;
        RECT 711.995 16.195 712.255 16.455 ;
        RECT 714.850 16.195 715.110 16.455 ;
        RECT 711.995 15.535 712.255 15.795 ;
        RECT 714.850 15.535 715.110 15.795 ;
        RECT 711.995 14.875 712.255 15.135 ;
        RECT 714.850 14.875 715.110 15.135 ;
        RECT 711.995 14.215 712.255 14.475 ;
        RECT 714.850 14.215 715.110 14.475 ;
        RECT 711.995 13.555 712.255 13.815 ;
        RECT 714.850 13.555 715.110 13.815 ;
        RECT 711.995 12.895 712.255 13.155 ;
        RECT 714.850 12.895 715.110 13.155 ;
        RECT 711.995 12.235 712.255 12.495 ;
        RECT 714.850 12.235 715.110 12.495 ;
        RECT 711.995 11.575 712.255 11.835 ;
        RECT 714.850 11.575 715.110 11.835 ;
        RECT 711.995 10.915 712.255 11.175 ;
        RECT 714.850 10.915 715.110 11.175 ;
        RECT 711.995 10.255 712.255 10.515 ;
        RECT 714.850 10.255 715.110 10.515 ;
        RECT 711.995 9.595 712.255 9.855 ;
        RECT 714.850 9.595 715.110 9.855 ;
        RECT 711.995 8.935 712.255 9.195 ;
        RECT 714.850 8.935 715.110 9.195 ;
        RECT 716.635 55.175 716.895 55.435 ;
        RECT 716.635 54.515 716.895 54.775 ;
        RECT 716.635 53.855 716.895 54.115 ;
        RECT 716.635 53.195 716.895 53.455 ;
        RECT 716.635 52.535 716.895 52.795 ;
        RECT 716.635 51.875 716.895 52.135 ;
        RECT 716.635 51.215 716.895 51.475 ;
        RECT 716.635 50.555 716.895 50.815 ;
        RECT 715.610 39.765 715.870 40.025 ;
        RECT 715.610 39.105 715.870 39.365 ;
        RECT 715.610 38.445 715.870 38.705 ;
        RECT 716.635 18.175 716.895 18.435 ;
        RECT 716.635 17.515 716.895 17.775 ;
        RECT 716.635 16.855 716.895 17.115 ;
        RECT 716.635 16.195 716.895 16.455 ;
        RECT 716.635 15.535 716.895 15.795 ;
        RECT 716.635 14.875 716.895 15.135 ;
        RECT 716.635 14.215 716.895 14.475 ;
        RECT 716.635 13.555 716.895 13.815 ;
        RECT 716.635 12.895 716.895 13.155 ;
        RECT 716.635 12.235 716.895 12.495 ;
        RECT 716.635 11.575 716.895 11.835 ;
        RECT 716.635 10.915 716.895 11.175 ;
        RECT 716.635 10.255 716.895 10.515 ;
        RECT 716.635 9.595 716.895 9.855 ;
        RECT 716.635 8.935 716.895 9.195 ;
        RECT 4.670 8.150 4.930 8.410 ;
        RECT 4.670 7.490 4.930 7.750 ;
        RECT 4.670 6.830 4.930 7.090 ;
        RECT 0.910 4.750 1.170 5.010 ;
        RECT 2.050 4.750 2.310 5.010 ;
        RECT 3.545 4.160 3.805 4.420 ;
        RECT 22.860 8.150 23.120 8.410 ;
        RECT 22.860 7.490 23.120 7.750 ;
        RECT 22.860 6.830 23.120 7.090 ;
        RECT 8.090 4.780 8.350 5.040 ;
        RECT 8.750 4.780 9.010 5.040 ;
        RECT 9.410 4.780 9.670 5.040 ;
        RECT 14.620 4.750 14.880 5.010 ;
        RECT 15.280 4.750 15.540 5.010 ;
        RECT 15.940 4.750 16.200 5.010 ;
        RECT 17.980 4.750 18.240 5.010 ;
        RECT 18.640 4.750 18.900 5.010 ;
        RECT 19.300 4.750 19.560 5.010 ;
        RECT 4.230 3.480 4.490 3.740 ;
        RECT 4.640 2.820 4.900 3.080 ;
        RECT 7.115 3.005 7.375 3.265 ;
        RECT 9.905 2.995 10.165 3.255 ;
        RECT 3.875 2.005 4.135 2.265 ;
        RECT 0.910 0.830 1.170 1.090 ;
        RECT 2.050 0.830 2.310 1.090 ;
        RECT 7.685 2.295 7.945 2.555 ;
        RECT 11.590 2.830 12.890 3.090 ;
        RECT 15.005 2.830 15.265 3.090 ;
        RECT 12.150 1.590 12.410 1.850 ;
        RECT 16.780 1.830 17.040 2.090 ;
        RECT 20.090 3.830 20.350 4.090 ;
        RECT 21.735 4.160 21.995 4.420 ;
        RECT 38.810 8.150 39.070 8.410 ;
        RECT 38.810 7.490 39.070 7.750 ;
        RECT 38.810 6.830 39.070 7.090 ;
        RECT 26.280 4.780 26.540 5.040 ;
        RECT 26.940 4.780 27.200 5.040 ;
        RECT 27.600 4.780 27.860 5.040 ;
        RECT 32.810 4.750 33.070 5.010 ;
        RECT 33.470 4.750 33.730 5.010 ;
        RECT 34.130 4.750 34.390 5.010 ;
        RECT 36.190 4.750 36.450 5.010 ;
        RECT 22.420 3.480 22.680 3.740 ;
        RECT 18.365 2.830 18.625 3.090 ;
        RECT 22.830 2.820 23.090 3.080 ;
        RECT 25.305 3.005 25.565 3.265 ;
        RECT 28.095 2.995 28.355 3.255 ;
        RECT 22.065 2.005 22.325 2.265 ;
        RECT 7.490 0.830 7.750 1.090 ;
        RECT 8.150 0.830 8.410 1.090 ;
        RECT 8.810 0.830 9.070 1.090 ;
        RECT 14.360 0.830 14.620 1.090 ;
        RECT 15.680 0.830 15.940 1.090 ;
        RECT 17.720 0.830 17.980 1.090 ;
        RECT 19.040 0.830 19.300 1.090 ;
        RECT 25.875 2.295 26.135 2.555 ;
        RECT 29.780 2.830 31.080 3.090 ;
        RECT 37.685 4.160 37.945 4.420 ;
        RECT 53.640 8.150 53.900 8.410 ;
        RECT 53.640 7.490 53.900 7.750 ;
        RECT 53.640 6.830 53.900 7.090 ;
        RECT 42.230 4.780 42.490 5.040 ;
        RECT 42.890 4.780 43.150 5.040 ;
        RECT 43.550 4.780 43.810 5.040 ;
        RECT 48.760 4.750 49.020 5.010 ;
        RECT 49.420 4.750 49.680 5.010 ;
        RECT 50.080 4.750 50.340 5.010 ;
        RECT 38.370 3.480 38.630 3.740 ;
        RECT 33.195 2.830 33.455 3.090 ;
        RECT 30.340 1.590 30.600 1.850 ;
        RECT 34.970 1.830 35.230 2.090 ;
        RECT 38.780 2.820 39.040 3.080 ;
        RECT 41.255 3.005 41.515 3.265 ;
        RECT 44.045 2.995 44.305 3.255 ;
        RECT 38.015 2.005 38.275 2.265 ;
        RECT 25.680 0.830 25.940 1.090 ;
        RECT 26.340 0.830 26.600 1.090 ;
        RECT 27.000 0.830 27.260 1.090 ;
        RECT 32.550 0.830 32.810 1.090 ;
        RECT 33.870 0.830 34.130 1.090 ;
        RECT 36.190 0.830 36.450 1.090 ;
        RECT 41.825 2.295 42.085 2.555 ;
        RECT 45.730 2.830 47.030 3.090 ;
        RECT 52.515 4.160 52.775 4.420 ;
        RECT 72.950 8.150 73.210 8.410 ;
        RECT 72.950 7.490 73.210 7.750 ;
        RECT 72.950 6.830 73.210 7.090 ;
        RECT 57.060 4.780 57.320 5.040 ;
        RECT 57.720 4.780 57.980 5.040 ;
        RECT 58.380 4.780 58.640 5.040 ;
        RECT 63.590 4.750 63.850 5.010 ;
        RECT 64.250 4.750 64.510 5.010 ;
        RECT 64.910 4.750 65.170 5.010 ;
        RECT 66.950 4.750 67.210 5.010 ;
        RECT 67.610 4.750 67.870 5.010 ;
        RECT 68.270 4.750 68.530 5.010 ;
        RECT 70.330 4.750 70.590 5.010 ;
        RECT 53.200 3.480 53.460 3.740 ;
        RECT 49.145 2.830 49.405 3.090 ;
        RECT 53.610 2.820 53.870 3.080 ;
        RECT 56.085 3.005 56.345 3.265 ;
        RECT 58.875 2.995 59.135 3.255 ;
        RECT 46.290 1.590 46.550 1.850 ;
        RECT 50.920 1.830 51.180 2.090 ;
        RECT 52.845 2.005 53.105 2.265 ;
        RECT 41.630 0.830 41.890 1.090 ;
        RECT 42.290 0.830 42.550 1.090 ;
        RECT 42.950 0.830 43.210 1.090 ;
        RECT 48.500 0.830 48.760 1.090 ;
        RECT 49.820 0.830 50.080 1.090 ;
        RECT 56.655 2.295 56.915 2.555 ;
        RECT 60.560 2.830 61.860 3.090 ;
        RECT 63.975 2.830 64.235 3.090 ;
        RECT 61.120 1.590 61.380 1.850 ;
        RECT 65.750 1.830 66.010 2.090 ;
        RECT 69.060 3.830 69.320 4.090 ;
        RECT 71.825 4.160 72.085 4.420 ;
        RECT 87.780 8.150 88.040 8.410 ;
        RECT 87.780 7.490 88.040 7.750 ;
        RECT 87.780 6.830 88.040 7.090 ;
        RECT 76.370 4.780 76.630 5.040 ;
        RECT 77.030 4.780 77.290 5.040 ;
        RECT 77.690 4.780 77.950 5.040 ;
        RECT 82.900 4.750 83.160 5.010 ;
        RECT 83.560 4.750 83.820 5.010 ;
        RECT 84.220 4.750 84.480 5.010 ;
        RECT 72.510 3.480 72.770 3.740 ;
        RECT 67.335 2.830 67.595 3.090 ;
        RECT 72.920 2.820 73.180 3.080 ;
        RECT 75.395 3.005 75.655 3.265 ;
        RECT 78.185 2.995 78.445 3.255 ;
        RECT 72.155 2.005 72.415 2.265 ;
        RECT 56.460 0.830 56.720 1.090 ;
        RECT 57.120 0.830 57.380 1.090 ;
        RECT 57.780 0.830 58.040 1.090 ;
        RECT 63.330 0.830 63.590 1.090 ;
        RECT 64.650 0.830 64.910 1.090 ;
        RECT 66.690 0.830 66.950 1.090 ;
        RECT 68.010 0.830 68.270 1.090 ;
        RECT 70.330 0.830 70.590 1.090 ;
        RECT 75.965 2.295 76.225 2.555 ;
        RECT 79.870 2.830 81.170 3.090 ;
        RECT 86.655 4.160 86.915 4.420 ;
        RECT 107.090 8.150 107.350 8.410 ;
        RECT 107.090 7.490 107.350 7.750 ;
        RECT 107.090 6.830 107.350 7.090 ;
        RECT 91.200 4.780 91.460 5.040 ;
        RECT 91.860 4.780 92.120 5.040 ;
        RECT 92.520 4.780 92.780 5.040 ;
        RECT 97.730 4.750 97.990 5.010 ;
        RECT 98.390 4.750 98.650 5.010 ;
        RECT 99.050 4.750 99.310 5.010 ;
        RECT 101.090 4.750 101.350 5.010 ;
        RECT 101.750 4.750 102.010 5.010 ;
        RECT 102.410 4.750 102.670 5.010 ;
        RECT 104.470 4.750 104.730 5.010 ;
        RECT 87.340 3.480 87.600 3.740 ;
        RECT 83.285 2.830 83.545 3.090 ;
        RECT 87.750 2.820 88.010 3.080 ;
        RECT 90.225 3.005 90.485 3.265 ;
        RECT 93.015 2.995 93.275 3.255 ;
        RECT 80.430 1.590 80.690 1.850 ;
        RECT 85.060 1.830 85.320 2.090 ;
        RECT 86.985 2.005 87.245 2.265 ;
        RECT 75.770 0.830 76.030 1.090 ;
        RECT 76.430 0.830 76.690 1.090 ;
        RECT 77.090 0.830 77.350 1.090 ;
        RECT 82.640 0.830 82.900 1.090 ;
        RECT 83.960 0.830 84.220 1.090 ;
        RECT 90.795 2.295 91.055 2.555 ;
        RECT 94.700 2.830 96.000 3.090 ;
        RECT 98.115 2.830 98.375 3.090 ;
        RECT 95.260 1.590 95.520 1.850 ;
        RECT 99.890 1.830 100.150 2.090 ;
        RECT 103.200 3.830 103.460 4.090 ;
        RECT 105.965 4.160 106.225 4.420 ;
        RECT 121.920 8.150 122.180 8.410 ;
        RECT 121.920 7.490 122.180 7.750 ;
        RECT 121.920 6.830 122.180 7.090 ;
        RECT 110.510 4.780 110.770 5.040 ;
        RECT 111.170 4.780 111.430 5.040 ;
        RECT 111.830 4.780 112.090 5.040 ;
        RECT 117.040 4.750 117.300 5.010 ;
        RECT 117.700 4.750 117.960 5.010 ;
        RECT 118.360 4.750 118.620 5.010 ;
        RECT 106.650 3.480 106.910 3.740 ;
        RECT 101.475 2.830 101.735 3.090 ;
        RECT 107.060 2.820 107.320 3.080 ;
        RECT 109.535 3.005 109.795 3.265 ;
        RECT 112.325 2.995 112.585 3.255 ;
        RECT 106.295 2.005 106.555 2.265 ;
        RECT 90.600 0.830 90.860 1.090 ;
        RECT 91.260 0.830 91.520 1.090 ;
        RECT 91.920 0.830 92.180 1.090 ;
        RECT 97.470 0.830 97.730 1.090 ;
        RECT 98.790 0.830 99.050 1.090 ;
        RECT 100.830 0.830 101.090 1.090 ;
        RECT 102.150 0.830 102.410 1.090 ;
        RECT 104.470 0.830 104.730 1.090 ;
        RECT 110.105 2.295 110.365 2.555 ;
        RECT 114.010 2.830 115.310 3.090 ;
        RECT 120.795 4.160 121.055 4.420 ;
        RECT 125.340 4.780 125.600 5.040 ;
        RECT 126.000 4.780 126.260 5.040 ;
        RECT 126.660 4.780 126.920 5.040 ;
        RECT 131.870 4.750 132.130 5.010 ;
        RECT 132.530 4.750 132.790 5.010 ;
        RECT 133.190 4.750 133.450 5.010 ;
        RECT 135.250 4.750 135.510 5.010 ;
        RECT 136.250 4.750 136.510 5.010 ;
        RECT 136.910 4.750 137.170 5.010 ;
        RECT 137.570 4.750 137.830 5.010 ;
        RECT 138.490 4.750 138.750 5.010 ;
        RECT 139.150 4.750 139.410 5.010 ;
        RECT 139.810 4.750 140.070 5.010 ;
        RECT 140.830 4.750 141.090 5.010 ;
        RECT 141.490 4.750 141.750 5.010 ;
        RECT 142.150 4.750 142.410 5.010 ;
        RECT 144.090 4.750 144.350 5.010 ;
        RECT 144.750 4.750 145.010 5.010 ;
        RECT 145.410 4.750 145.670 5.010 ;
        RECT 146.330 4.750 146.590 5.010 ;
        RECT 146.990 4.750 147.250 5.010 ;
        RECT 147.650 4.750 147.910 5.010 ;
        RECT 148.570 4.750 148.830 5.010 ;
        RECT 149.230 4.750 149.490 5.010 ;
        RECT 149.890 4.750 150.150 5.010 ;
        RECT 150.810 4.750 151.070 5.010 ;
        RECT 151.470 4.750 151.730 5.010 ;
        RECT 152.130 4.750 152.390 5.010 ;
        RECT 153.050 4.750 153.310 5.010 ;
        RECT 153.710 4.750 153.970 5.010 ;
        RECT 154.370 4.750 154.630 5.010 ;
        RECT 155.410 4.750 155.670 5.010 ;
        RECT 156.410 4.750 156.670 5.010 ;
        RECT 157.070 4.750 157.330 5.010 ;
        RECT 157.730 4.750 157.990 5.010 ;
        RECT 158.650 4.750 158.910 5.010 ;
        RECT 159.310 4.750 159.570 5.010 ;
        RECT 159.970 4.750 160.230 5.010 ;
        RECT 160.890 4.750 161.150 5.010 ;
        RECT 161.550 4.750 161.810 5.010 ;
        RECT 162.210 4.750 162.470 5.010 ;
        RECT 163.130 4.750 163.390 5.010 ;
        RECT 163.790 4.750 164.050 5.010 ;
        RECT 164.450 4.750 164.710 5.010 ;
        RECT 165.370 4.750 165.630 5.010 ;
        RECT 166.030 4.750 166.290 5.010 ;
        RECT 166.690 4.750 166.950 5.010 ;
        RECT 167.610 4.750 167.870 5.010 ;
        RECT 168.270 4.750 168.530 5.010 ;
        RECT 168.930 4.750 169.190 5.010 ;
        RECT 169.850 4.750 170.110 5.010 ;
        RECT 170.510 4.750 170.770 5.010 ;
        RECT 171.170 4.750 171.430 5.010 ;
        RECT 172.090 4.750 172.350 5.010 ;
        RECT 172.750 4.750 173.010 5.010 ;
        RECT 173.410 4.750 173.670 5.010 ;
        RECT 174.330 4.750 174.590 5.010 ;
        RECT 174.990 4.750 175.250 5.010 ;
        RECT 175.650 4.750 175.910 5.010 ;
        RECT 176.690 4.750 176.950 5.010 ;
        RECT 177.690 4.750 177.950 5.010 ;
        RECT 178.350 4.750 178.610 5.010 ;
        RECT 179.010 4.750 179.270 5.010 ;
        RECT 179.930 4.750 180.190 5.010 ;
        RECT 180.590 4.750 180.850 5.010 ;
        RECT 181.250 4.750 181.510 5.010 ;
        RECT 182.270 4.750 182.530 5.010 ;
        RECT 182.930 4.750 183.190 5.010 ;
        RECT 183.590 4.750 183.850 5.010 ;
        RECT 185.530 4.750 185.790 5.010 ;
        RECT 186.190 4.750 186.450 5.010 ;
        RECT 186.850 4.750 187.110 5.010 ;
        RECT 187.770 4.750 188.030 5.010 ;
        RECT 188.430 4.750 188.690 5.010 ;
        RECT 189.090 4.750 189.350 5.010 ;
        RECT 190.010 4.750 190.270 5.010 ;
        RECT 190.670 4.750 190.930 5.010 ;
        RECT 191.330 4.750 191.590 5.010 ;
        RECT 192.250 4.750 192.510 5.010 ;
        RECT 192.910 4.750 193.170 5.010 ;
        RECT 193.570 4.750 193.830 5.010 ;
        RECT 194.490 4.750 194.750 5.010 ;
        RECT 195.150 4.750 195.410 5.010 ;
        RECT 195.810 4.750 196.070 5.010 ;
        RECT 196.850 4.750 197.110 5.010 ;
        RECT 197.850 4.750 198.110 5.010 ;
        RECT 198.510 4.750 198.770 5.010 ;
        RECT 199.170 4.750 199.430 5.010 ;
        RECT 200.090 4.750 200.350 5.010 ;
        RECT 200.750 4.750 201.010 5.010 ;
        RECT 201.410 4.750 201.670 5.010 ;
        RECT 202.330 4.750 202.590 5.010 ;
        RECT 202.990 4.750 203.250 5.010 ;
        RECT 203.650 4.750 203.910 5.010 ;
        RECT 204.570 4.750 204.830 5.010 ;
        RECT 205.230 4.750 205.490 5.010 ;
        RECT 205.890 4.750 206.150 5.010 ;
        RECT 206.810 4.750 207.070 5.010 ;
        RECT 207.470 4.750 207.730 5.010 ;
        RECT 208.130 4.750 208.390 5.010 ;
        RECT 209.050 4.750 209.310 5.010 ;
        RECT 209.710 4.750 209.970 5.010 ;
        RECT 210.370 4.750 210.630 5.010 ;
        RECT 211.290 4.750 211.550 5.010 ;
        RECT 211.950 4.750 212.210 5.010 ;
        RECT 212.610 4.750 212.870 5.010 ;
        RECT 213.530 4.750 213.790 5.010 ;
        RECT 214.190 4.750 214.450 5.010 ;
        RECT 214.850 4.750 215.110 5.010 ;
        RECT 215.770 4.750 216.030 5.010 ;
        RECT 216.430 4.750 216.690 5.010 ;
        RECT 217.090 4.750 217.350 5.010 ;
        RECT 218.130 4.750 218.390 5.010 ;
        RECT 219.130 4.750 219.390 5.010 ;
        RECT 219.790 4.750 220.050 5.010 ;
        RECT 220.450 4.750 220.710 5.010 ;
        RECT 221.370 4.750 221.630 5.010 ;
        RECT 222.030 4.750 222.290 5.010 ;
        RECT 222.690 4.750 222.950 5.010 ;
        RECT 223.610 4.750 223.870 5.010 ;
        RECT 224.270 4.750 224.530 5.010 ;
        RECT 224.930 4.750 225.190 5.010 ;
        RECT 225.950 4.750 226.210 5.010 ;
        RECT 226.610 4.750 226.870 5.010 ;
        RECT 227.270 4.750 227.530 5.010 ;
        RECT 229.210 4.750 229.470 5.010 ;
        RECT 229.870 4.750 230.130 5.010 ;
        RECT 230.530 4.750 230.790 5.010 ;
        RECT 231.450 4.750 231.710 5.010 ;
        RECT 232.110 4.750 232.370 5.010 ;
        RECT 232.770 4.750 233.030 5.010 ;
        RECT 233.690 4.750 233.950 5.010 ;
        RECT 234.350 4.750 234.610 5.010 ;
        RECT 235.010 4.750 235.270 5.010 ;
        RECT 235.930 4.750 236.190 5.010 ;
        RECT 236.590 4.750 236.850 5.010 ;
        RECT 237.250 4.750 237.510 5.010 ;
        RECT 238.290 4.750 238.550 5.010 ;
        RECT 239.290 4.750 239.550 5.010 ;
        RECT 239.950 4.750 240.210 5.010 ;
        RECT 240.610 4.750 240.870 5.010 ;
        RECT 241.530 4.750 241.790 5.010 ;
        RECT 242.190 4.750 242.450 5.010 ;
        RECT 242.850 4.750 243.110 5.010 ;
        RECT 243.770 4.750 244.030 5.010 ;
        RECT 244.430 4.750 244.690 5.010 ;
        RECT 245.090 4.750 245.350 5.010 ;
        RECT 246.010 4.750 246.270 5.010 ;
        RECT 246.670 4.750 246.930 5.010 ;
        RECT 247.330 4.750 247.590 5.010 ;
        RECT 248.250 4.750 248.510 5.010 ;
        RECT 248.910 4.750 249.170 5.010 ;
        RECT 249.570 4.750 249.830 5.010 ;
        RECT 250.490 4.750 250.750 5.010 ;
        RECT 251.150 4.750 251.410 5.010 ;
        RECT 251.810 4.750 252.070 5.010 ;
        RECT 252.730 4.750 252.990 5.010 ;
        RECT 253.390 4.750 253.650 5.010 ;
        RECT 254.050 4.750 254.310 5.010 ;
        RECT 254.970 4.750 255.230 5.010 ;
        RECT 255.630 4.750 255.890 5.010 ;
        RECT 256.290 4.750 256.550 5.010 ;
        RECT 257.210 4.750 257.470 5.010 ;
        RECT 257.870 4.750 258.130 5.010 ;
        RECT 258.530 4.750 258.790 5.010 ;
        RECT 259.570 4.750 259.830 5.010 ;
        RECT 260.570 4.750 260.830 5.010 ;
        RECT 261.230 4.750 261.490 5.010 ;
        RECT 261.890 4.750 262.150 5.010 ;
        RECT 262.810 4.750 263.070 5.010 ;
        RECT 263.470 4.750 263.730 5.010 ;
        RECT 264.130 4.750 264.390 5.010 ;
        RECT 265.050 4.750 265.310 5.010 ;
        RECT 265.710 4.750 265.970 5.010 ;
        RECT 266.370 4.750 266.630 5.010 ;
        RECT 267.390 4.750 267.650 5.010 ;
        RECT 268.050 4.750 268.310 5.010 ;
        RECT 268.710 4.750 268.970 5.010 ;
        RECT 270.650 4.750 270.910 5.010 ;
        RECT 271.310 4.750 271.570 5.010 ;
        RECT 271.970 4.750 272.230 5.010 ;
        RECT 272.890 4.750 273.150 5.010 ;
        RECT 273.550 4.750 273.810 5.010 ;
        RECT 274.210 4.750 274.470 5.010 ;
        RECT 275.130 4.750 275.390 5.010 ;
        RECT 275.790 4.750 276.050 5.010 ;
        RECT 276.450 4.750 276.710 5.010 ;
        RECT 277.370 4.750 277.630 5.010 ;
        RECT 278.030 4.750 278.290 5.010 ;
        RECT 278.690 4.750 278.950 5.010 ;
        RECT 279.730 4.750 279.990 5.010 ;
        RECT 280.730 4.750 280.990 5.010 ;
        RECT 281.390 4.750 281.650 5.010 ;
        RECT 282.050 4.750 282.310 5.010 ;
        RECT 282.970 4.750 283.230 5.010 ;
        RECT 283.630 4.750 283.890 5.010 ;
        RECT 284.290 4.750 284.550 5.010 ;
        RECT 285.210 4.750 285.470 5.010 ;
        RECT 285.870 4.750 286.130 5.010 ;
        RECT 286.530 4.750 286.790 5.010 ;
        RECT 287.450 4.750 287.710 5.010 ;
        RECT 288.110 4.750 288.370 5.010 ;
        RECT 288.770 4.750 289.030 5.010 ;
        RECT 289.690 4.750 289.950 5.010 ;
        RECT 290.350 4.750 290.610 5.010 ;
        RECT 291.010 4.750 291.270 5.010 ;
        RECT 291.930 4.750 292.190 5.010 ;
        RECT 292.590 4.750 292.850 5.010 ;
        RECT 293.250 4.750 293.510 5.010 ;
        RECT 294.170 4.750 294.430 5.010 ;
        RECT 294.830 4.750 295.090 5.010 ;
        RECT 295.490 4.750 295.750 5.010 ;
        RECT 296.410 4.750 296.670 5.010 ;
        RECT 297.070 4.750 297.330 5.010 ;
        RECT 297.730 4.750 297.990 5.010 ;
        RECT 298.650 4.750 298.910 5.010 ;
        RECT 299.310 4.750 299.570 5.010 ;
        RECT 299.970 4.750 300.230 5.010 ;
        RECT 301.010 4.750 301.270 5.010 ;
        RECT 302.010 4.750 302.270 5.010 ;
        RECT 302.670 4.750 302.930 5.010 ;
        RECT 303.330 4.750 303.590 5.010 ;
        RECT 304.250 4.750 304.510 5.010 ;
        RECT 304.910 4.750 305.170 5.010 ;
        RECT 305.570 4.750 305.830 5.010 ;
        RECT 306.490 4.750 306.750 5.010 ;
        RECT 307.150 4.750 307.410 5.010 ;
        RECT 307.810 4.750 308.070 5.010 ;
        RECT 308.730 4.750 308.990 5.010 ;
        RECT 309.390 4.750 309.650 5.010 ;
        RECT 310.050 4.750 310.310 5.010 ;
        RECT 311.070 4.750 311.330 5.010 ;
        RECT 311.730 4.750 311.990 5.010 ;
        RECT 312.390 4.750 312.650 5.010 ;
        RECT 314.330 4.750 314.590 5.010 ;
        RECT 314.990 4.750 315.250 5.010 ;
        RECT 315.650 4.750 315.910 5.010 ;
        RECT 316.570 4.750 316.830 5.010 ;
        RECT 317.230 4.750 317.490 5.010 ;
        RECT 317.890 4.750 318.150 5.010 ;
        RECT 318.810 4.750 319.070 5.010 ;
        RECT 319.470 4.750 319.730 5.010 ;
        RECT 320.130 4.750 320.390 5.010 ;
        RECT 321.170 4.750 321.430 5.010 ;
        RECT 322.170 4.750 322.430 5.010 ;
        RECT 322.830 4.750 323.090 5.010 ;
        RECT 323.490 4.750 323.750 5.010 ;
        RECT 324.410 4.750 324.670 5.010 ;
        RECT 325.070 4.750 325.330 5.010 ;
        RECT 325.730 4.750 325.990 5.010 ;
        RECT 326.650 4.750 326.910 5.010 ;
        RECT 327.310 4.750 327.570 5.010 ;
        RECT 327.970 4.750 328.230 5.010 ;
        RECT 328.890 4.750 329.150 5.010 ;
        RECT 329.550 4.750 329.810 5.010 ;
        RECT 330.210 4.750 330.470 5.010 ;
        RECT 331.130 4.750 331.390 5.010 ;
        RECT 331.790 4.750 332.050 5.010 ;
        RECT 332.450 4.750 332.710 5.010 ;
        RECT 333.370 4.750 333.630 5.010 ;
        RECT 334.030 4.750 334.290 5.010 ;
        RECT 334.690 4.750 334.950 5.010 ;
        RECT 335.610 4.750 335.870 5.010 ;
        RECT 336.270 4.750 336.530 5.010 ;
        RECT 336.930 4.750 337.190 5.010 ;
        RECT 337.850 4.750 338.110 5.010 ;
        RECT 338.510 4.750 338.770 5.010 ;
        RECT 339.170 4.750 339.430 5.010 ;
        RECT 340.090 4.750 340.350 5.010 ;
        RECT 340.750 4.750 341.010 5.010 ;
        RECT 341.410 4.750 341.670 5.010 ;
        RECT 342.450 4.750 342.710 5.010 ;
        RECT 343.450 4.750 343.710 5.010 ;
        RECT 344.110 4.750 344.370 5.010 ;
        RECT 344.770 4.750 345.030 5.010 ;
        RECT 345.690 4.750 345.950 5.010 ;
        RECT 346.350 4.750 346.610 5.010 ;
        RECT 347.010 4.750 347.270 5.010 ;
        RECT 347.930 4.750 348.190 5.010 ;
        RECT 348.590 4.750 348.850 5.010 ;
        RECT 349.250 4.750 349.510 5.010 ;
        RECT 350.170 4.750 350.430 5.010 ;
        RECT 350.830 4.750 351.090 5.010 ;
        RECT 351.490 4.750 351.750 5.010 ;
        RECT 352.510 4.750 352.770 5.010 ;
        RECT 353.170 4.750 353.430 5.010 ;
        RECT 353.830 4.750 354.090 5.010 ;
        RECT 355.770 4.750 356.030 5.010 ;
        RECT 356.430 4.750 356.690 5.010 ;
        RECT 357.090 4.750 357.350 5.010 ;
        RECT 358.010 4.750 358.270 5.010 ;
        RECT 358.670 4.750 358.930 5.010 ;
        RECT 359.330 4.750 359.590 5.010 ;
        RECT 360.250 4.750 360.510 5.010 ;
        RECT 360.910 4.750 361.170 5.010 ;
        RECT 361.570 4.750 361.830 5.010 ;
        RECT 362.610 4.750 362.870 5.010 ;
        RECT 363.610 4.750 363.870 5.010 ;
        RECT 364.270 4.750 364.530 5.010 ;
        RECT 364.930 4.750 365.190 5.010 ;
        RECT 365.850 4.750 366.110 5.010 ;
        RECT 366.510 4.750 366.770 5.010 ;
        RECT 367.170 4.750 367.430 5.010 ;
        RECT 368.090 4.750 368.350 5.010 ;
        RECT 368.750 4.750 369.010 5.010 ;
        RECT 369.410 4.750 369.670 5.010 ;
        RECT 370.330 4.750 370.590 5.010 ;
        RECT 370.990 4.750 371.250 5.010 ;
        RECT 371.650 4.750 371.910 5.010 ;
        RECT 372.570 4.750 372.830 5.010 ;
        RECT 373.230 4.750 373.490 5.010 ;
        RECT 373.890 4.750 374.150 5.010 ;
        RECT 374.810 4.750 375.070 5.010 ;
        RECT 375.470 4.750 375.730 5.010 ;
        RECT 376.130 4.750 376.390 5.010 ;
        RECT 377.050 4.750 377.310 5.010 ;
        RECT 377.710 4.750 377.970 5.010 ;
        RECT 378.370 4.750 378.630 5.010 ;
        RECT 379.290 4.750 379.550 5.010 ;
        RECT 379.950 4.750 380.210 5.010 ;
        RECT 380.610 4.750 380.870 5.010 ;
        RECT 381.530 4.750 381.790 5.010 ;
        RECT 382.190 4.750 382.450 5.010 ;
        RECT 382.850 4.750 383.110 5.010 ;
        RECT 383.890 4.750 384.150 5.010 ;
        RECT 384.890 4.750 385.150 5.010 ;
        RECT 385.550 4.750 385.810 5.010 ;
        RECT 386.210 4.750 386.470 5.010 ;
        RECT 387.130 4.750 387.390 5.010 ;
        RECT 387.790 4.750 388.050 5.010 ;
        RECT 388.450 4.750 388.710 5.010 ;
        RECT 389.370 4.750 389.630 5.010 ;
        RECT 390.030 4.750 390.290 5.010 ;
        RECT 390.690 4.750 390.950 5.010 ;
        RECT 391.610 4.750 391.870 5.010 ;
        RECT 392.270 4.750 392.530 5.010 ;
        RECT 392.930 4.750 393.190 5.010 ;
        RECT 393.850 4.750 394.110 5.010 ;
        RECT 394.510 4.750 394.770 5.010 ;
        RECT 395.170 4.750 395.430 5.010 ;
        RECT 396.190 4.750 396.450 5.010 ;
        RECT 396.850 4.750 397.110 5.010 ;
        RECT 397.510 4.750 397.770 5.010 ;
        RECT 399.450 4.750 399.710 5.010 ;
        RECT 400.110 4.750 400.370 5.010 ;
        RECT 400.770 4.750 401.030 5.010 ;
        RECT 401.690 4.750 401.950 5.010 ;
        RECT 402.350 4.750 402.610 5.010 ;
        RECT 403.010 4.750 403.270 5.010 ;
        RECT 404.050 4.750 404.310 5.010 ;
        RECT 405.050 4.750 405.310 5.010 ;
        RECT 405.710 4.750 405.970 5.010 ;
        RECT 406.370 4.750 406.630 5.010 ;
        RECT 407.290 4.750 407.550 5.010 ;
        RECT 407.950 4.750 408.210 5.010 ;
        RECT 408.610 4.750 408.870 5.010 ;
        RECT 409.530 4.750 409.790 5.010 ;
        RECT 410.190 4.750 410.450 5.010 ;
        RECT 410.850 4.750 411.110 5.010 ;
        RECT 411.770 4.750 412.030 5.010 ;
        RECT 412.430 4.750 412.690 5.010 ;
        RECT 413.090 4.750 413.350 5.010 ;
        RECT 414.010 4.750 414.270 5.010 ;
        RECT 414.670 4.750 414.930 5.010 ;
        RECT 415.330 4.750 415.590 5.010 ;
        RECT 416.250 4.750 416.510 5.010 ;
        RECT 416.910 4.750 417.170 5.010 ;
        RECT 417.570 4.750 417.830 5.010 ;
        RECT 418.490 4.750 418.750 5.010 ;
        RECT 419.150 4.750 419.410 5.010 ;
        RECT 419.810 4.750 420.070 5.010 ;
        RECT 420.730 4.750 420.990 5.010 ;
        RECT 421.390 4.750 421.650 5.010 ;
        RECT 422.050 4.750 422.310 5.010 ;
        RECT 422.970 4.750 423.230 5.010 ;
        RECT 423.630 4.750 423.890 5.010 ;
        RECT 424.290 4.750 424.550 5.010 ;
        RECT 425.330 4.750 425.590 5.010 ;
        RECT 426.330 4.750 426.590 5.010 ;
        RECT 426.990 4.750 427.250 5.010 ;
        RECT 427.650 4.750 427.910 5.010 ;
        RECT 428.570 4.750 428.830 5.010 ;
        RECT 429.230 4.750 429.490 5.010 ;
        RECT 429.890 4.750 430.150 5.010 ;
        RECT 430.810 4.750 431.070 5.010 ;
        RECT 431.470 4.750 431.730 5.010 ;
        RECT 432.130 4.750 432.390 5.010 ;
        RECT 433.050 4.750 433.310 5.010 ;
        RECT 433.710 4.750 433.970 5.010 ;
        RECT 434.370 4.750 434.630 5.010 ;
        RECT 435.290 4.750 435.550 5.010 ;
        RECT 435.950 4.750 436.210 5.010 ;
        RECT 436.610 4.750 436.870 5.010 ;
        RECT 437.630 4.750 437.890 5.010 ;
        RECT 438.290 4.750 438.550 5.010 ;
        RECT 438.950 4.750 439.210 5.010 ;
        RECT 440.890 4.750 441.150 5.010 ;
        RECT 441.550 4.750 441.810 5.010 ;
        RECT 442.210 4.750 442.470 5.010 ;
        RECT 443.130 4.750 443.390 5.010 ;
        RECT 443.790 4.750 444.050 5.010 ;
        RECT 444.450 4.750 444.710 5.010 ;
        RECT 445.490 4.750 445.750 5.010 ;
        RECT 446.490 4.750 446.750 5.010 ;
        RECT 447.150 4.750 447.410 5.010 ;
        RECT 447.810 4.750 448.070 5.010 ;
        RECT 448.730 4.750 448.990 5.010 ;
        RECT 449.390 4.750 449.650 5.010 ;
        RECT 450.050 4.750 450.310 5.010 ;
        RECT 450.970 4.750 451.230 5.010 ;
        RECT 451.630 4.750 451.890 5.010 ;
        RECT 452.290 4.750 452.550 5.010 ;
        RECT 453.210 4.750 453.470 5.010 ;
        RECT 453.870 4.750 454.130 5.010 ;
        RECT 454.530 4.750 454.790 5.010 ;
        RECT 455.450 4.750 455.710 5.010 ;
        RECT 456.110 4.750 456.370 5.010 ;
        RECT 456.770 4.750 457.030 5.010 ;
        RECT 457.690 4.750 457.950 5.010 ;
        RECT 458.350 4.750 458.610 5.010 ;
        RECT 459.010 4.750 459.270 5.010 ;
        RECT 459.930 4.750 460.190 5.010 ;
        RECT 460.590 4.750 460.850 5.010 ;
        RECT 461.250 4.750 461.510 5.010 ;
        RECT 462.170 4.750 462.430 5.010 ;
        RECT 462.830 4.750 463.090 5.010 ;
        RECT 463.490 4.750 463.750 5.010 ;
        RECT 464.410 4.750 464.670 5.010 ;
        RECT 465.070 4.750 465.330 5.010 ;
        RECT 465.730 4.750 465.990 5.010 ;
        RECT 466.770 4.750 467.030 5.010 ;
        RECT 467.770 4.750 468.030 5.010 ;
        RECT 468.430 4.750 468.690 5.010 ;
        RECT 469.090 4.750 469.350 5.010 ;
        RECT 470.010 4.750 470.270 5.010 ;
        RECT 470.670 4.750 470.930 5.010 ;
        RECT 471.330 4.750 471.590 5.010 ;
        RECT 472.250 4.750 472.510 5.010 ;
        RECT 472.910 4.750 473.170 5.010 ;
        RECT 473.570 4.750 473.830 5.010 ;
        RECT 474.490 4.750 474.750 5.010 ;
        RECT 475.150 4.750 475.410 5.010 ;
        RECT 475.810 4.750 476.070 5.010 ;
        RECT 476.730 4.750 476.990 5.010 ;
        RECT 477.390 4.750 477.650 5.010 ;
        RECT 478.050 4.750 478.310 5.010 ;
        RECT 478.970 4.750 479.230 5.010 ;
        RECT 479.630 4.750 479.890 5.010 ;
        RECT 480.290 4.750 480.550 5.010 ;
        RECT 481.310 4.750 481.570 5.010 ;
        RECT 481.970 4.750 482.230 5.010 ;
        RECT 482.630 4.750 482.890 5.010 ;
        RECT 484.570 4.750 484.830 5.010 ;
        RECT 485.230 4.750 485.490 5.010 ;
        RECT 485.890 4.750 486.150 5.010 ;
        RECT 486.930 4.750 487.190 5.010 ;
        RECT 487.930 4.750 488.190 5.010 ;
        RECT 488.590 4.750 488.850 5.010 ;
        RECT 489.250 4.750 489.510 5.010 ;
        RECT 490.170 4.750 490.430 5.010 ;
        RECT 490.830 4.750 491.090 5.010 ;
        RECT 491.490 4.750 491.750 5.010 ;
        RECT 492.410 4.750 492.670 5.010 ;
        RECT 493.070 4.750 493.330 5.010 ;
        RECT 493.730 4.750 493.990 5.010 ;
        RECT 494.650 4.750 494.910 5.010 ;
        RECT 495.310 4.750 495.570 5.010 ;
        RECT 495.970 4.750 496.230 5.010 ;
        RECT 496.890 4.750 497.150 5.010 ;
        RECT 497.550 4.750 497.810 5.010 ;
        RECT 498.210 4.750 498.470 5.010 ;
        RECT 499.130 4.750 499.390 5.010 ;
        RECT 499.790 4.750 500.050 5.010 ;
        RECT 500.450 4.750 500.710 5.010 ;
        RECT 501.370 4.750 501.630 5.010 ;
        RECT 502.030 4.750 502.290 5.010 ;
        RECT 502.690 4.750 502.950 5.010 ;
        RECT 503.610 4.750 503.870 5.010 ;
        RECT 504.270 4.750 504.530 5.010 ;
        RECT 504.930 4.750 505.190 5.010 ;
        RECT 505.850 4.750 506.110 5.010 ;
        RECT 506.510 4.750 506.770 5.010 ;
        RECT 507.170 4.750 507.430 5.010 ;
        RECT 508.210 4.750 508.470 5.010 ;
        RECT 509.210 4.750 509.470 5.010 ;
        RECT 509.870 4.750 510.130 5.010 ;
        RECT 510.530 4.750 510.790 5.010 ;
        RECT 511.450 4.750 511.710 5.010 ;
        RECT 512.110 4.750 512.370 5.010 ;
        RECT 512.770 4.750 513.030 5.010 ;
        RECT 513.690 4.750 513.950 5.010 ;
        RECT 514.350 4.750 514.610 5.010 ;
        RECT 515.010 4.750 515.270 5.010 ;
        RECT 515.930 4.750 516.190 5.010 ;
        RECT 516.590 4.750 516.850 5.010 ;
        RECT 517.250 4.750 517.510 5.010 ;
        RECT 518.170 4.750 518.430 5.010 ;
        RECT 518.830 4.750 519.090 5.010 ;
        RECT 519.490 4.750 519.750 5.010 ;
        RECT 520.410 4.750 520.670 5.010 ;
        RECT 521.070 4.750 521.330 5.010 ;
        RECT 521.730 4.750 521.990 5.010 ;
        RECT 522.750 4.750 523.010 5.010 ;
        RECT 523.410 4.750 523.670 5.010 ;
        RECT 524.070 4.750 524.330 5.010 ;
        RECT 526.010 4.750 526.270 5.010 ;
        RECT 526.670 4.750 526.930 5.010 ;
        RECT 527.330 4.750 527.590 5.010 ;
        RECT 528.370 4.750 528.630 5.010 ;
        RECT 529.370 4.750 529.630 5.010 ;
        RECT 530.030 4.750 530.290 5.010 ;
        RECT 530.690 4.750 530.950 5.010 ;
        RECT 531.610 4.750 531.870 5.010 ;
        RECT 532.270 4.750 532.530 5.010 ;
        RECT 532.930 4.750 533.190 5.010 ;
        RECT 533.850 4.750 534.110 5.010 ;
        RECT 534.510 4.750 534.770 5.010 ;
        RECT 535.170 4.750 535.430 5.010 ;
        RECT 536.090 4.750 536.350 5.010 ;
        RECT 536.750 4.750 537.010 5.010 ;
        RECT 537.410 4.750 537.670 5.010 ;
        RECT 538.330 4.750 538.590 5.010 ;
        RECT 538.990 4.750 539.250 5.010 ;
        RECT 539.650 4.750 539.910 5.010 ;
        RECT 540.570 4.750 540.830 5.010 ;
        RECT 541.230 4.750 541.490 5.010 ;
        RECT 541.890 4.750 542.150 5.010 ;
        RECT 542.810 4.750 543.070 5.010 ;
        RECT 543.470 4.750 543.730 5.010 ;
        RECT 544.130 4.750 544.390 5.010 ;
        RECT 545.050 4.750 545.310 5.010 ;
        RECT 545.710 4.750 545.970 5.010 ;
        RECT 546.370 4.750 546.630 5.010 ;
        RECT 547.290 4.750 547.550 5.010 ;
        RECT 547.950 4.750 548.210 5.010 ;
        RECT 548.610 4.750 548.870 5.010 ;
        RECT 549.650 4.750 549.910 5.010 ;
        RECT 550.650 4.750 550.910 5.010 ;
        RECT 551.310 4.750 551.570 5.010 ;
        RECT 551.970 4.750 552.230 5.010 ;
        RECT 552.890 4.750 553.150 5.010 ;
        RECT 553.550 4.750 553.810 5.010 ;
        RECT 554.210 4.750 554.470 5.010 ;
        RECT 555.130 4.750 555.390 5.010 ;
        RECT 555.790 4.750 556.050 5.010 ;
        RECT 556.450 4.750 556.710 5.010 ;
        RECT 557.370 4.750 557.630 5.010 ;
        RECT 558.030 4.750 558.290 5.010 ;
        RECT 558.690 4.750 558.950 5.010 ;
        RECT 559.610 4.750 559.870 5.010 ;
        RECT 560.270 4.750 560.530 5.010 ;
        RECT 560.930 4.750 561.190 5.010 ;
        RECT 561.850 4.750 562.110 5.010 ;
        RECT 562.510 4.750 562.770 5.010 ;
        RECT 563.170 4.750 563.430 5.010 ;
        RECT 564.090 4.750 564.350 5.010 ;
        RECT 564.750 4.750 565.010 5.010 ;
        RECT 565.410 4.750 565.670 5.010 ;
        RECT 566.430 4.750 566.690 5.010 ;
        RECT 567.090 4.750 567.350 5.010 ;
        RECT 567.750 4.750 568.010 5.010 ;
        RECT 569.810 4.750 570.070 5.010 ;
        RECT 570.810 4.750 571.070 5.010 ;
        RECT 571.470 4.750 571.730 5.010 ;
        RECT 572.130 4.750 572.390 5.010 ;
        RECT 573.050 4.750 573.310 5.010 ;
        RECT 573.710 4.750 573.970 5.010 ;
        RECT 574.370 4.750 574.630 5.010 ;
        RECT 575.290 4.750 575.550 5.010 ;
        RECT 575.950 4.750 576.210 5.010 ;
        RECT 576.610 4.750 576.870 5.010 ;
        RECT 577.530 4.750 577.790 5.010 ;
        RECT 578.190 4.750 578.450 5.010 ;
        RECT 578.850 4.750 579.110 5.010 ;
        RECT 579.770 4.750 580.030 5.010 ;
        RECT 580.430 4.750 580.690 5.010 ;
        RECT 581.090 4.750 581.350 5.010 ;
        RECT 582.010 4.750 582.270 5.010 ;
        RECT 582.670 4.750 582.930 5.010 ;
        RECT 583.330 4.750 583.590 5.010 ;
        RECT 584.250 4.750 584.510 5.010 ;
        RECT 584.910 4.750 585.170 5.010 ;
        RECT 585.570 4.750 585.830 5.010 ;
        RECT 586.490 4.750 586.750 5.010 ;
        RECT 587.150 4.750 587.410 5.010 ;
        RECT 587.810 4.750 588.070 5.010 ;
        RECT 588.730 4.750 588.990 5.010 ;
        RECT 589.390 4.750 589.650 5.010 ;
        RECT 590.050 4.750 590.310 5.010 ;
        RECT 591.090 4.750 591.350 5.010 ;
        RECT 592.090 4.750 592.350 5.010 ;
        RECT 592.750 4.750 593.010 5.010 ;
        RECT 593.410 4.750 593.670 5.010 ;
        RECT 594.330 4.750 594.590 5.010 ;
        RECT 594.990 4.750 595.250 5.010 ;
        RECT 595.650 4.750 595.910 5.010 ;
        RECT 596.570 4.750 596.830 5.010 ;
        RECT 597.230 4.750 597.490 5.010 ;
        RECT 597.890 4.750 598.150 5.010 ;
        RECT 598.810 4.750 599.070 5.010 ;
        RECT 599.470 4.750 599.730 5.010 ;
        RECT 600.130 4.750 600.390 5.010 ;
        RECT 601.050 4.750 601.310 5.010 ;
        RECT 601.710 4.750 601.970 5.010 ;
        RECT 602.370 4.750 602.630 5.010 ;
        RECT 603.290 4.750 603.550 5.010 ;
        RECT 603.950 4.750 604.210 5.010 ;
        RECT 604.610 4.750 604.870 5.010 ;
        RECT 605.530 4.750 605.790 5.010 ;
        RECT 606.190 4.750 606.450 5.010 ;
        RECT 606.850 4.750 607.110 5.010 ;
        RECT 607.870 4.750 608.130 5.010 ;
        RECT 608.530 4.750 608.790 5.010 ;
        RECT 609.190 4.750 609.450 5.010 ;
        RECT 611.250 4.750 611.510 5.010 ;
        RECT 612.250 4.750 612.510 5.010 ;
        RECT 612.910 4.750 613.170 5.010 ;
        RECT 613.570 4.750 613.830 5.010 ;
        RECT 614.490 4.750 614.750 5.010 ;
        RECT 615.150 4.750 615.410 5.010 ;
        RECT 615.810 4.750 616.070 5.010 ;
        RECT 616.730 4.750 616.990 5.010 ;
        RECT 617.390 4.750 617.650 5.010 ;
        RECT 618.050 4.750 618.310 5.010 ;
        RECT 618.970 4.750 619.230 5.010 ;
        RECT 619.630 4.750 619.890 5.010 ;
        RECT 620.290 4.750 620.550 5.010 ;
        RECT 621.210 4.750 621.470 5.010 ;
        RECT 621.870 4.750 622.130 5.010 ;
        RECT 622.530 4.750 622.790 5.010 ;
        RECT 623.450 4.750 623.710 5.010 ;
        RECT 624.110 4.750 624.370 5.010 ;
        RECT 624.770 4.750 625.030 5.010 ;
        RECT 625.690 4.750 625.950 5.010 ;
        RECT 626.350 4.750 626.610 5.010 ;
        RECT 627.010 4.750 627.270 5.010 ;
        RECT 627.930 4.750 628.190 5.010 ;
        RECT 628.590 4.750 628.850 5.010 ;
        RECT 629.250 4.750 629.510 5.010 ;
        RECT 630.170 4.750 630.430 5.010 ;
        RECT 630.830 4.750 631.090 5.010 ;
        RECT 631.490 4.750 631.750 5.010 ;
        RECT 632.530 4.750 632.790 5.010 ;
        RECT 633.530 4.750 633.790 5.010 ;
        RECT 634.190 4.750 634.450 5.010 ;
        RECT 634.850 4.750 635.110 5.010 ;
        RECT 635.770 4.750 636.030 5.010 ;
        RECT 636.430 4.750 636.690 5.010 ;
        RECT 637.090 4.750 637.350 5.010 ;
        RECT 638.010 4.750 638.270 5.010 ;
        RECT 638.670 4.750 638.930 5.010 ;
        RECT 639.330 4.750 639.590 5.010 ;
        RECT 640.250 4.750 640.510 5.010 ;
        RECT 640.910 4.750 641.170 5.010 ;
        RECT 641.570 4.750 641.830 5.010 ;
        RECT 642.490 4.750 642.750 5.010 ;
        RECT 643.150 4.750 643.410 5.010 ;
        RECT 643.810 4.750 644.070 5.010 ;
        RECT 644.730 4.750 644.990 5.010 ;
        RECT 645.390 4.750 645.650 5.010 ;
        RECT 646.050 4.750 646.310 5.010 ;
        RECT 646.970 4.750 647.230 5.010 ;
        RECT 647.630 4.750 647.890 5.010 ;
        RECT 648.290 4.750 648.550 5.010 ;
        RECT 649.210 4.750 649.470 5.010 ;
        RECT 649.870 4.750 650.130 5.010 ;
        RECT 650.530 4.750 650.790 5.010 ;
        RECT 651.550 4.750 651.810 5.010 ;
        RECT 652.210 4.750 652.470 5.010 ;
        RECT 652.870 4.750 653.130 5.010 ;
        RECT 654.930 4.750 655.190 5.010 ;
        RECT 655.930 4.750 656.190 5.010 ;
        RECT 656.590 4.750 656.850 5.010 ;
        RECT 657.250 4.750 657.510 5.010 ;
        RECT 658.170 4.750 658.430 5.010 ;
        RECT 658.830 4.750 659.090 5.010 ;
        RECT 659.490 4.750 659.750 5.010 ;
        RECT 660.410 4.750 660.670 5.010 ;
        RECT 661.070 4.750 661.330 5.010 ;
        RECT 661.730 4.750 661.990 5.010 ;
        RECT 662.650 4.750 662.910 5.010 ;
        RECT 663.310 4.750 663.570 5.010 ;
        RECT 663.970 4.750 664.230 5.010 ;
        RECT 664.890 4.750 665.150 5.010 ;
        RECT 665.550 4.750 665.810 5.010 ;
        RECT 666.210 4.750 666.470 5.010 ;
        RECT 667.130 4.750 667.390 5.010 ;
        RECT 667.790 4.750 668.050 5.010 ;
        RECT 668.450 4.750 668.710 5.010 ;
        RECT 669.370 4.750 669.630 5.010 ;
        RECT 670.030 4.750 670.290 5.010 ;
        RECT 670.690 4.750 670.950 5.010 ;
        RECT 671.610 4.750 671.870 5.010 ;
        RECT 672.270 4.750 672.530 5.010 ;
        RECT 672.930 4.750 673.190 5.010 ;
        RECT 673.850 4.750 674.110 5.010 ;
        RECT 674.510 4.750 674.770 5.010 ;
        RECT 675.170 4.750 675.430 5.010 ;
        RECT 676.210 4.750 676.470 5.010 ;
        RECT 677.210 4.750 677.470 5.010 ;
        RECT 677.870 4.750 678.130 5.010 ;
        RECT 678.530 4.750 678.790 5.010 ;
        RECT 679.550 4.750 679.810 5.010 ;
        RECT 121.480 3.480 121.740 3.740 ;
        RECT 117.425 2.830 117.685 3.090 ;
        RECT 121.890 2.820 122.150 3.080 ;
        RECT 124.365 3.005 124.625 3.265 ;
        RECT 127.155 2.995 127.415 3.255 ;
        RECT 114.570 1.590 114.830 1.850 ;
        RECT 119.200 1.830 119.460 2.090 ;
        RECT 121.125 2.005 121.385 2.265 ;
        RECT 109.910 0.830 110.170 1.090 ;
        RECT 110.570 0.830 110.830 1.090 ;
        RECT 111.230 0.830 111.490 1.090 ;
        RECT 116.780 0.830 117.040 1.090 ;
        RECT 118.100 0.830 118.360 1.090 ;
        RECT 124.935 2.295 125.195 2.555 ;
        RECT 128.840 2.830 130.140 3.090 ;
        RECT 132.255 2.830 132.515 3.090 ;
        RECT 129.400 1.590 129.660 1.850 ;
        RECT 134.030 1.830 134.290 2.090 ;
        RECT 142.940 3.830 143.200 4.090 ;
        RECT 141.215 2.830 141.475 3.090 ;
        RECT 184.380 3.830 184.640 4.090 ;
        RECT 182.655 2.830 182.915 3.090 ;
        RECT 228.060 3.830 228.320 4.090 ;
        RECT 226.335 2.830 226.595 3.090 ;
        RECT 269.500 3.830 269.760 4.090 ;
        RECT 267.775 2.830 268.035 3.090 ;
        RECT 313.180 3.830 313.440 4.090 ;
        RECT 311.455 2.830 311.715 3.090 ;
        RECT 354.620 3.830 354.880 4.090 ;
        RECT 352.895 2.830 353.155 3.090 ;
        RECT 398.300 3.830 398.560 4.090 ;
        RECT 396.575 2.830 396.835 3.090 ;
        RECT 439.740 3.830 440.000 4.090 ;
        RECT 438.015 2.830 438.275 3.090 ;
        RECT 483.420 3.830 483.680 4.090 ;
        RECT 481.695 2.830 481.955 3.090 ;
        RECT 524.860 3.830 525.120 4.090 ;
        RECT 523.135 2.830 523.395 3.090 ;
        RECT 568.540 3.830 568.800 4.090 ;
        RECT 566.815 2.830 567.075 3.090 ;
        RECT 609.980 3.830 610.240 4.090 ;
        RECT 608.255 2.830 608.515 3.090 ;
        RECT 653.660 3.830 653.920 4.090 ;
        RECT 651.935 2.830 652.195 3.090 ;
        RECT 124.740 0.830 125.000 1.090 ;
        RECT 125.400 0.830 125.660 1.090 ;
        RECT 126.060 0.830 126.320 1.090 ;
        RECT 131.610 0.830 131.870 1.090 ;
        RECT 132.930 0.830 133.190 1.090 ;
        RECT 135.250 0.830 135.510 1.090 ;
        RECT 136.250 0.830 136.510 1.090 ;
        RECT 136.910 0.830 137.170 1.090 ;
        RECT 137.570 0.830 137.830 1.090 ;
        RECT 138.490 0.830 138.750 1.090 ;
        RECT 139.150 0.830 139.410 1.090 ;
        RECT 139.810 0.830 140.070 1.090 ;
        RECT 140.570 0.830 140.830 1.090 ;
        RECT 141.890 0.830 142.150 1.090 ;
        RECT 144.090 0.830 144.350 1.090 ;
        RECT 144.750 0.830 145.010 1.090 ;
        RECT 145.410 0.830 145.670 1.090 ;
        RECT 146.330 0.830 146.590 1.090 ;
        RECT 146.990 0.830 147.250 1.090 ;
        RECT 147.650 0.830 147.910 1.090 ;
        RECT 148.570 0.830 148.830 1.090 ;
        RECT 149.230 0.830 149.490 1.090 ;
        RECT 149.890 0.830 150.150 1.090 ;
        RECT 150.810 0.830 151.070 1.090 ;
        RECT 151.470 0.830 151.730 1.090 ;
        RECT 152.130 0.830 152.390 1.090 ;
        RECT 153.050 0.830 153.310 1.090 ;
        RECT 153.710 0.830 153.970 1.090 ;
        RECT 154.370 0.830 154.630 1.090 ;
        RECT 155.410 0.830 155.670 1.090 ;
        RECT 156.410 0.830 156.670 1.090 ;
        RECT 157.070 0.830 157.330 1.090 ;
        RECT 157.730 0.830 157.990 1.090 ;
        RECT 158.650 0.830 158.910 1.090 ;
        RECT 159.310 0.830 159.570 1.090 ;
        RECT 159.970 0.830 160.230 1.090 ;
        RECT 160.890 0.830 161.150 1.090 ;
        RECT 161.550 0.830 161.810 1.090 ;
        RECT 162.210 0.830 162.470 1.090 ;
        RECT 163.130 0.830 163.390 1.090 ;
        RECT 163.790 0.830 164.050 1.090 ;
        RECT 164.450 0.830 164.710 1.090 ;
        RECT 165.370 0.830 165.630 1.090 ;
        RECT 166.030 0.830 166.290 1.090 ;
        RECT 166.690 0.830 166.950 1.090 ;
        RECT 167.610 0.830 167.870 1.090 ;
        RECT 168.270 0.830 168.530 1.090 ;
        RECT 168.930 0.830 169.190 1.090 ;
        RECT 169.850 0.830 170.110 1.090 ;
        RECT 170.510 0.830 170.770 1.090 ;
        RECT 171.170 0.830 171.430 1.090 ;
        RECT 172.090 0.830 172.350 1.090 ;
        RECT 172.750 0.830 173.010 1.090 ;
        RECT 173.410 0.830 173.670 1.090 ;
        RECT 174.330 0.830 174.590 1.090 ;
        RECT 174.990 0.830 175.250 1.090 ;
        RECT 175.650 0.830 175.910 1.090 ;
        RECT 176.690 0.830 176.950 1.090 ;
        RECT 177.690 0.830 177.950 1.090 ;
        RECT 178.350 0.830 178.610 1.090 ;
        RECT 179.010 0.830 179.270 1.090 ;
        RECT 179.930 0.830 180.190 1.090 ;
        RECT 180.590 0.830 180.850 1.090 ;
        RECT 181.250 0.830 181.510 1.090 ;
        RECT 182.010 0.830 182.270 1.090 ;
        RECT 183.330 0.830 183.590 1.090 ;
        RECT 185.530 0.830 185.790 1.090 ;
        RECT 186.190 0.830 186.450 1.090 ;
        RECT 186.850 0.830 187.110 1.090 ;
        RECT 187.770 0.830 188.030 1.090 ;
        RECT 188.430 0.830 188.690 1.090 ;
        RECT 189.090 0.830 189.350 1.090 ;
        RECT 190.010 0.830 190.270 1.090 ;
        RECT 190.670 0.830 190.930 1.090 ;
        RECT 191.330 0.830 191.590 1.090 ;
        RECT 192.250 0.830 192.510 1.090 ;
        RECT 192.910 0.830 193.170 1.090 ;
        RECT 193.570 0.830 193.830 1.090 ;
        RECT 194.490 0.830 194.750 1.090 ;
        RECT 195.150 0.830 195.410 1.090 ;
        RECT 195.810 0.830 196.070 1.090 ;
        RECT 196.850 0.830 197.110 1.090 ;
        RECT 197.850 0.830 198.110 1.090 ;
        RECT 198.510 0.830 198.770 1.090 ;
        RECT 199.170 0.830 199.430 1.090 ;
        RECT 200.090 0.830 200.350 1.090 ;
        RECT 200.750 0.830 201.010 1.090 ;
        RECT 201.410 0.830 201.670 1.090 ;
        RECT 202.330 0.830 202.590 1.090 ;
        RECT 202.990 0.830 203.250 1.090 ;
        RECT 203.650 0.830 203.910 1.090 ;
        RECT 204.570 0.830 204.830 1.090 ;
        RECT 205.230 0.830 205.490 1.090 ;
        RECT 205.890 0.830 206.150 1.090 ;
        RECT 206.810 0.830 207.070 1.090 ;
        RECT 207.470 0.830 207.730 1.090 ;
        RECT 208.130 0.830 208.390 1.090 ;
        RECT 209.050 0.830 209.310 1.090 ;
        RECT 209.710 0.830 209.970 1.090 ;
        RECT 210.370 0.830 210.630 1.090 ;
        RECT 211.290 0.830 211.550 1.090 ;
        RECT 211.950 0.830 212.210 1.090 ;
        RECT 212.610 0.830 212.870 1.090 ;
        RECT 213.530 0.830 213.790 1.090 ;
        RECT 214.190 0.830 214.450 1.090 ;
        RECT 214.850 0.830 215.110 1.090 ;
        RECT 215.770 0.830 216.030 1.090 ;
        RECT 216.430 0.830 216.690 1.090 ;
        RECT 217.090 0.830 217.350 1.090 ;
        RECT 218.130 0.830 218.390 1.090 ;
        RECT 219.130 0.830 219.390 1.090 ;
        RECT 219.790 0.830 220.050 1.090 ;
        RECT 220.450 0.830 220.710 1.090 ;
        RECT 221.370 0.830 221.630 1.090 ;
        RECT 222.030 0.830 222.290 1.090 ;
        RECT 222.690 0.830 222.950 1.090 ;
        RECT 223.610 0.830 223.870 1.090 ;
        RECT 224.270 0.830 224.530 1.090 ;
        RECT 224.930 0.830 225.190 1.090 ;
        RECT 225.690 0.830 225.950 1.090 ;
        RECT 227.010 0.830 227.270 1.090 ;
        RECT 229.210 0.830 229.470 1.090 ;
        RECT 229.870 0.830 230.130 1.090 ;
        RECT 230.530 0.830 230.790 1.090 ;
        RECT 231.450 0.830 231.710 1.090 ;
        RECT 232.110 0.830 232.370 1.090 ;
        RECT 232.770 0.830 233.030 1.090 ;
        RECT 233.690 0.830 233.950 1.090 ;
        RECT 234.350 0.830 234.610 1.090 ;
        RECT 235.010 0.830 235.270 1.090 ;
        RECT 235.930 0.830 236.190 1.090 ;
        RECT 236.590 0.830 236.850 1.090 ;
        RECT 237.250 0.830 237.510 1.090 ;
        RECT 238.290 0.830 238.550 1.090 ;
        RECT 239.290 0.830 239.550 1.090 ;
        RECT 239.950 0.830 240.210 1.090 ;
        RECT 240.610 0.830 240.870 1.090 ;
        RECT 241.530 0.830 241.790 1.090 ;
        RECT 242.190 0.830 242.450 1.090 ;
        RECT 242.850 0.830 243.110 1.090 ;
        RECT 243.770 0.830 244.030 1.090 ;
        RECT 244.430 0.830 244.690 1.090 ;
        RECT 245.090 0.830 245.350 1.090 ;
        RECT 246.010 0.830 246.270 1.090 ;
        RECT 246.670 0.830 246.930 1.090 ;
        RECT 247.330 0.830 247.590 1.090 ;
        RECT 248.250 0.830 248.510 1.090 ;
        RECT 248.910 0.830 249.170 1.090 ;
        RECT 249.570 0.830 249.830 1.090 ;
        RECT 250.490 0.830 250.750 1.090 ;
        RECT 251.150 0.830 251.410 1.090 ;
        RECT 251.810 0.830 252.070 1.090 ;
        RECT 252.730 0.830 252.990 1.090 ;
        RECT 253.390 0.830 253.650 1.090 ;
        RECT 254.050 0.830 254.310 1.090 ;
        RECT 254.970 0.830 255.230 1.090 ;
        RECT 255.630 0.830 255.890 1.090 ;
        RECT 256.290 0.830 256.550 1.090 ;
        RECT 257.210 0.830 257.470 1.090 ;
        RECT 257.870 0.830 258.130 1.090 ;
        RECT 258.530 0.830 258.790 1.090 ;
        RECT 259.570 0.830 259.830 1.090 ;
        RECT 260.570 0.830 260.830 1.090 ;
        RECT 261.230 0.830 261.490 1.090 ;
        RECT 261.890 0.830 262.150 1.090 ;
        RECT 262.810 0.830 263.070 1.090 ;
        RECT 263.470 0.830 263.730 1.090 ;
        RECT 264.130 0.830 264.390 1.090 ;
        RECT 265.050 0.830 265.310 1.090 ;
        RECT 265.710 0.830 265.970 1.090 ;
        RECT 266.370 0.830 266.630 1.090 ;
        RECT 267.130 0.830 267.390 1.090 ;
        RECT 268.450 0.830 268.710 1.090 ;
        RECT 270.650 0.830 270.910 1.090 ;
        RECT 271.310 0.830 271.570 1.090 ;
        RECT 271.970 0.830 272.230 1.090 ;
        RECT 272.890 0.830 273.150 1.090 ;
        RECT 273.550 0.830 273.810 1.090 ;
        RECT 274.210 0.830 274.470 1.090 ;
        RECT 275.130 0.830 275.390 1.090 ;
        RECT 275.790 0.830 276.050 1.090 ;
        RECT 276.450 0.830 276.710 1.090 ;
        RECT 277.370 0.830 277.630 1.090 ;
        RECT 278.030 0.830 278.290 1.090 ;
        RECT 278.690 0.830 278.950 1.090 ;
        RECT 279.730 0.830 279.990 1.090 ;
        RECT 280.730 0.830 280.990 1.090 ;
        RECT 281.390 0.830 281.650 1.090 ;
        RECT 282.050 0.830 282.310 1.090 ;
        RECT 282.970 0.830 283.230 1.090 ;
        RECT 283.630 0.830 283.890 1.090 ;
        RECT 284.290 0.830 284.550 1.090 ;
        RECT 285.210 0.830 285.470 1.090 ;
        RECT 285.870 0.830 286.130 1.090 ;
        RECT 286.530 0.830 286.790 1.090 ;
        RECT 287.450 0.830 287.710 1.090 ;
        RECT 288.110 0.830 288.370 1.090 ;
        RECT 288.770 0.830 289.030 1.090 ;
        RECT 289.690 0.830 289.950 1.090 ;
        RECT 290.350 0.830 290.610 1.090 ;
        RECT 291.010 0.830 291.270 1.090 ;
        RECT 291.930 0.830 292.190 1.090 ;
        RECT 292.590 0.830 292.850 1.090 ;
        RECT 293.250 0.830 293.510 1.090 ;
        RECT 294.170 0.830 294.430 1.090 ;
        RECT 294.830 0.830 295.090 1.090 ;
        RECT 295.490 0.830 295.750 1.090 ;
        RECT 296.410 0.830 296.670 1.090 ;
        RECT 297.070 0.830 297.330 1.090 ;
        RECT 297.730 0.830 297.990 1.090 ;
        RECT 298.650 0.830 298.910 1.090 ;
        RECT 299.310 0.830 299.570 1.090 ;
        RECT 299.970 0.830 300.230 1.090 ;
        RECT 301.010 0.830 301.270 1.090 ;
        RECT 302.010 0.830 302.270 1.090 ;
        RECT 302.670 0.830 302.930 1.090 ;
        RECT 303.330 0.830 303.590 1.090 ;
        RECT 304.250 0.830 304.510 1.090 ;
        RECT 304.910 0.830 305.170 1.090 ;
        RECT 305.570 0.830 305.830 1.090 ;
        RECT 306.490 0.830 306.750 1.090 ;
        RECT 307.150 0.830 307.410 1.090 ;
        RECT 307.810 0.830 308.070 1.090 ;
        RECT 308.730 0.830 308.990 1.090 ;
        RECT 309.390 0.830 309.650 1.090 ;
        RECT 310.050 0.830 310.310 1.090 ;
        RECT 310.810 0.830 311.070 1.090 ;
        RECT 312.130 0.830 312.390 1.090 ;
        RECT 314.330 0.830 314.590 1.090 ;
        RECT 314.990 0.830 315.250 1.090 ;
        RECT 315.650 0.830 315.910 1.090 ;
        RECT 316.570 0.830 316.830 1.090 ;
        RECT 317.230 0.830 317.490 1.090 ;
        RECT 317.890 0.830 318.150 1.090 ;
        RECT 318.810 0.830 319.070 1.090 ;
        RECT 319.470 0.830 319.730 1.090 ;
        RECT 320.130 0.830 320.390 1.090 ;
        RECT 321.170 0.830 321.430 1.090 ;
        RECT 322.170 0.830 322.430 1.090 ;
        RECT 322.830 0.830 323.090 1.090 ;
        RECT 323.490 0.830 323.750 1.090 ;
        RECT 324.410 0.830 324.670 1.090 ;
        RECT 325.070 0.830 325.330 1.090 ;
        RECT 325.730 0.830 325.990 1.090 ;
        RECT 326.650 0.830 326.910 1.090 ;
        RECT 327.310 0.830 327.570 1.090 ;
        RECT 327.970 0.830 328.230 1.090 ;
        RECT 328.890 0.830 329.150 1.090 ;
        RECT 329.550 0.830 329.810 1.090 ;
        RECT 330.210 0.830 330.470 1.090 ;
        RECT 331.130 0.830 331.390 1.090 ;
        RECT 331.790 0.830 332.050 1.090 ;
        RECT 332.450 0.830 332.710 1.090 ;
        RECT 333.370 0.830 333.630 1.090 ;
        RECT 334.030 0.830 334.290 1.090 ;
        RECT 334.690 0.830 334.950 1.090 ;
        RECT 335.610 0.830 335.870 1.090 ;
        RECT 336.270 0.830 336.530 1.090 ;
        RECT 336.930 0.830 337.190 1.090 ;
        RECT 337.850 0.830 338.110 1.090 ;
        RECT 338.510 0.830 338.770 1.090 ;
        RECT 339.170 0.830 339.430 1.090 ;
        RECT 340.090 0.830 340.350 1.090 ;
        RECT 340.750 0.830 341.010 1.090 ;
        RECT 341.410 0.830 341.670 1.090 ;
        RECT 342.450 0.830 342.710 1.090 ;
        RECT 343.450 0.830 343.710 1.090 ;
        RECT 344.110 0.830 344.370 1.090 ;
        RECT 344.770 0.830 345.030 1.090 ;
        RECT 345.690 0.830 345.950 1.090 ;
        RECT 346.350 0.830 346.610 1.090 ;
        RECT 347.010 0.830 347.270 1.090 ;
        RECT 347.930 0.830 348.190 1.090 ;
        RECT 348.590 0.830 348.850 1.090 ;
        RECT 349.250 0.830 349.510 1.090 ;
        RECT 350.170 0.830 350.430 1.090 ;
        RECT 350.830 0.830 351.090 1.090 ;
        RECT 351.490 0.830 351.750 1.090 ;
        RECT 352.250 0.830 352.510 1.090 ;
        RECT 353.570 0.830 353.830 1.090 ;
        RECT 355.770 0.830 356.030 1.090 ;
        RECT 356.430 0.830 356.690 1.090 ;
        RECT 357.090 0.830 357.350 1.090 ;
        RECT 358.010 0.830 358.270 1.090 ;
        RECT 358.670 0.830 358.930 1.090 ;
        RECT 359.330 0.830 359.590 1.090 ;
        RECT 360.250 0.830 360.510 1.090 ;
        RECT 360.910 0.830 361.170 1.090 ;
        RECT 361.570 0.830 361.830 1.090 ;
        RECT 362.610 0.830 362.870 1.090 ;
        RECT 363.610 0.830 363.870 1.090 ;
        RECT 364.270 0.830 364.530 1.090 ;
        RECT 364.930 0.830 365.190 1.090 ;
        RECT 365.850 0.830 366.110 1.090 ;
        RECT 366.510 0.830 366.770 1.090 ;
        RECT 367.170 0.830 367.430 1.090 ;
        RECT 368.090 0.830 368.350 1.090 ;
        RECT 368.750 0.830 369.010 1.090 ;
        RECT 369.410 0.830 369.670 1.090 ;
        RECT 370.330 0.830 370.590 1.090 ;
        RECT 370.990 0.830 371.250 1.090 ;
        RECT 371.650 0.830 371.910 1.090 ;
        RECT 372.570 0.830 372.830 1.090 ;
        RECT 373.230 0.830 373.490 1.090 ;
        RECT 373.890 0.830 374.150 1.090 ;
        RECT 374.810 0.830 375.070 1.090 ;
        RECT 375.470 0.830 375.730 1.090 ;
        RECT 376.130 0.830 376.390 1.090 ;
        RECT 377.050 0.830 377.310 1.090 ;
        RECT 377.710 0.830 377.970 1.090 ;
        RECT 378.370 0.830 378.630 1.090 ;
        RECT 379.290 0.830 379.550 1.090 ;
        RECT 379.950 0.830 380.210 1.090 ;
        RECT 380.610 0.830 380.870 1.090 ;
        RECT 381.530 0.830 381.790 1.090 ;
        RECT 382.190 0.830 382.450 1.090 ;
        RECT 382.850 0.830 383.110 1.090 ;
        RECT 383.890 0.830 384.150 1.090 ;
        RECT 384.890 0.830 385.150 1.090 ;
        RECT 385.550 0.830 385.810 1.090 ;
        RECT 386.210 0.830 386.470 1.090 ;
        RECT 387.130 0.830 387.390 1.090 ;
        RECT 387.790 0.830 388.050 1.090 ;
        RECT 388.450 0.830 388.710 1.090 ;
        RECT 389.370 0.830 389.630 1.090 ;
        RECT 390.030 0.830 390.290 1.090 ;
        RECT 390.690 0.830 390.950 1.090 ;
        RECT 391.610 0.830 391.870 1.090 ;
        RECT 392.270 0.830 392.530 1.090 ;
        RECT 392.930 0.830 393.190 1.090 ;
        RECT 393.850 0.830 394.110 1.090 ;
        RECT 394.510 0.830 394.770 1.090 ;
        RECT 395.170 0.830 395.430 1.090 ;
        RECT 395.930 0.830 396.190 1.090 ;
        RECT 397.250 0.830 397.510 1.090 ;
        RECT 399.450 0.830 399.710 1.090 ;
        RECT 400.110 0.830 400.370 1.090 ;
        RECT 400.770 0.830 401.030 1.090 ;
        RECT 401.690 0.830 401.950 1.090 ;
        RECT 402.350 0.830 402.610 1.090 ;
        RECT 403.010 0.830 403.270 1.090 ;
        RECT 404.050 0.830 404.310 1.090 ;
        RECT 405.050 0.830 405.310 1.090 ;
        RECT 405.710 0.830 405.970 1.090 ;
        RECT 406.370 0.830 406.630 1.090 ;
        RECT 407.290 0.830 407.550 1.090 ;
        RECT 407.950 0.830 408.210 1.090 ;
        RECT 408.610 0.830 408.870 1.090 ;
        RECT 409.530 0.830 409.790 1.090 ;
        RECT 410.190 0.830 410.450 1.090 ;
        RECT 410.850 0.830 411.110 1.090 ;
        RECT 411.770 0.830 412.030 1.090 ;
        RECT 412.430 0.830 412.690 1.090 ;
        RECT 413.090 0.830 413.350 1.090 ;
        RECT 414.010 0.830 414.270 1.090 ;
        RECT 414.670 0.830 414.930 1.090 ;
        RECT 415.330 0.830 415.590 1.090 ;
        RECT 416.250 0.830 416.510 1.090 ;
        RECT 416.910 0.830 417.170 1.090 ;
        RECT 417.570 0.830 417.830 1.090 ;
        RECT 418.490 0.830 418.750 1.090 ;
        RECT 419.150 0.830 419.410 1.090 ;
        RECT 419.810 0.830 420.070 1.090 ;
        RECT 420.730 0.830 420.990 1.090 ;
        RECT 421.390 0.830 421.650 1.090 ;
        RECT 422.050 0.830 422.310 1.090 ;
        RECT 422.970 0.830 423.230 1.090 ;
        RECT 423.630 0.830 423.890 1.090 ;
        RECT 424.290 0.830 424.550 1.090 ;
        RECT 425.330 0.830 425.590 1.090 ;
        RECT 426.330 0.830 426.590 1.090 ;
        RECT 426.990 0.830 427.250 1.090 ;
        RECT 427.650 0.830 427.910 1.090 ;
        RECT 428.570 0.830 428.830 1.090 ;
        RECT 429.230 0.830 429.490 1.090 ;
        RECT 429.890 0.830 430.150 1.090 ;
        RECT 430.810 0.830 431.070 1.090 ;
        RECT 431.470 0.830 431.730 1.090 ;
        RECT 432.130 0.830 432.390 1.090 ;
        RECT 433.050 0.830 433.310 1.090 ;
        RECT 433.710 0.830 433.970 1.090 ;
        RECT 434.370 0.830 434.630 1.090 ;
        RECT 435.290 0.830 435.550 1.090 ;
        RECT 435.950 0.830 436.210 1.090 ;
        RECT 436.610 0.830 436.870 1.090 ;
        RECT 437.370 0.830 437.630 1.090 ;
        RECT 438.690 0.830 438.950 1.090 ;
        RECT 440.890 0.830 441.150 1.090 ;
        RECT 441.550 0.830 441.810 1.090 ;
        RECT 442.210 0.830 442.470 1.090 ;
        RECT 443.130 0.830 443.390 1.090 ;
        RECT 443.790 0.830 444.050 1.090 ;
        RECT 444.450 0.830 444.710 1.090 ;
        RECT 445.490 0.830 445.750 1.090 ;
        RECT 446.490 0.830 446.750 1.090 ;
        RECT 447.150 0.830 447.410 1.090 ;
        RECT 447.810 0.830 448.070 1.090 ;
        RECT 448.730 0.830 448.990 1.090 ;
        RECT 449.390 0.830 449.650 1.090 ;
        RECT 450.050 0.830 450.310 1.090 ;
        RECT 450.970 0.830 451.230 1.090 ;
        RECT 451.630 0.830 451.890 1.090 ;
        RECT 452.290 0.830 452.550 1.090 ;
        RECT 453.210 0.830 453.470 1.090 ;
        RECT 453.870 0.830 454.130 1.090 ;
        RECT 454.530 0.830 454.790 1.090 ;
        RECT 455.450 0.830 455.710 1.090 ;
        RECT 456.110 0.830 456.370 1.090 ;
        RECT 456.770 0.830 457.030 1.090 ;
        RECT 457.690 0.830 457.950 1.090 ;
        RECT 458.350 0.830 458.610 1.090 ;
        RECT 459.010 0.830 459.270 1.090 ;
        RECT 459.930 0.830 460.190 1.090 ;
        RECT 460.590 0.830 460.850 1.090 ;
        RECT 461.250 0.830 461.510 1.090 ;
        RECT 462.170 0.830 462.430 1.090 ;
        RECT 462.830 0.830 463.090 1.090 ;
        RECT 463.490 0.830 463.750 1.090 ;
        RECT 464.410 0.830 464.670 1.090 ;
        RECT 465.070 0.830 465.330 1.090 ;
        RECT 465.730 0.830 465.990 1.090 ;
        RECT 466.770 0.830 467.030 1.090 ;
        RECT 467.770 0.830 468.030 1.090 ;
        RECT 468.430 0.830 468.690 1.090 ;
        RECT 469.090 0.830 469.350 1.090 ;
        RECT 470.010 0.830 470.270 1.090 ;
        RECT 470.670 0.830 470.930 1.090 ;
        RECT 471.330 0.830 471.590 1.090 ;
        RECT 472.250 0.830 472.510 1.090 ;
        RECT 472.910 0.830 473.170 1.090 ;
        RECT 473.570 0.830 473.830 1.090 ;
        RECT 474.490 0.830 474.750 1.090 ;
        RECT 475.150 0.830 475.410 1.090 ;
        RECT 475.810 0.830 476.070 1.090 ;
        RECT 476.730 0.830 476.990 1.090 ;
        RECT 477.390 0.830 477.650 1.090 ;
        RECT 478.050 0.830 478.310 1.090 ;
        RECT 478.970 0.830 479.230 1.090 ;
        RECT 479.630 0.830 479.890 1.090 ;
        RECT 480.290 0.830 480.550 1.090 ;
        RECT 481.050 0.830 481.310 1.090 ;
        RECT 482.370 0.830 482.630 1.090 ;
        RECT 484.570 0.830 484.830 1.090 ;
        RECT 485.230 0.830 485.490 1.090 ;
        RECT 485.890 0.830 486.150 1.090 ;
        RECT 486.930 0.830 487.190 1.090 ;
        RECT 487.930 0.830 488.190 1.090 ;
        RECT 488.590 0.830 488.850 1.090 ;
        RECT 489.250 0.830 489.510 1.090 ;
        RECT 490.170 0.830 490.430 1.090 ;
        RECT 490.830 0.830 491.090 1.090 ;
        RECT 491.490 0.830 491.750 1.090 ;
        RECT 492.410 0.830 492.670 1.090 ;
        RECT 493.070 0.830 493.330 1.090 ;
        RECT 493.730 0.830 493.990 1.090 ;
        RECT 494.650 0.830 494.910 1.090 ;
        RECT 495.310 0.830 495.570 1.090 ;
        RECT 495.970 0.830 496.230 1.090 ;
        RECT 496.890 0.830 497.150 1.090 ;
        RECT 497.550 0.830 497.810 1.090 ;
        RECT 498.210 0.830 498.470 1.090 ;
        RECT 499.130 0.830 499.390 1.090 ;
        RECT 499.790 0.830 500.050 1.090 ;
        RECT 500.450 0.830 500.710 1.090 ;
        RECT 501.370 0.830 501.630 1.090 ;
        RECT 502.030 0.830 502.290 1.090 ;
        RECT 502.690 0.830 502.950 1.090 ;
        RECT 503.610 0.830 503.870 1.090 ;
        RECT 504.270 0.830 504.530 1.090 ;
        RECT 504.930 0.830 505.190 1.090 ;
        RECT 505.850 0.830 506.110 1.090 ;
        RECT 506.510 0.830 506.770 1.090 ;
        RECT 507.170 0.830 507.430 1.090 ;
        RECT 508.210 0.830 508.470 1.090 ;
        RECT 509.210 0.830 509.470 1.090 ;
        RECT 509.870 0.830 510.130 1.090 ;
        RECT 510.530 0.830 510.790 1.090 ;
        RECT 511.450 0.830 511.710 1.090 ;
        RECT 512.110 0.830 512.370 1.090 ;
        RECT 512.770 0.830 513.030 1.090 ;
        RECT 513.690 0.830 513.950 1.090 ;
        RECT 514.350 0.830 514.610 1.090 ;
        RECT 515.010 0.830 515.270 1.090 ;
        RECT 515.930 0.830 516.190 1.090 ;
        RECT 516.590 0.830 516.850 1.090 ;
        RECT 517.250 0.830 517.510 1.090 ;
        RECT 518.170 0.830 518.430 1.090 ;
        RECT 518.830 0.830 519.090 1.090 ;
        RECT 519.490 0.830 519.750 1.090 ;
        RECT 520.410 0.830 520.670 1.090 ;
        RECT 521.070 0.830 521.330 1.090 ;
        RECT 521.730 0.830 521.990 1.090 ;
        RECT 522.490 0.830 522.750 1.090 ;
        RECT 523.810 0.830 524.070 1.090 ;
        RECT 526.010 0.830 526.270 1.090 ;
        RECT 526.670 0.830 526.930 1.090 ;
        RECT 527.330 0.830 527.590 1.090 ;
        RECT 528.370 0.830 528.630 1.090 ;
        RECT 529.370 0.830 529.630 1.090 ;
        RECT 530.030 0.830 530.290 1.090 ;
        RECT 530.690 0.830 530.950 1.090 ;
        RECT 531.610 0.830 531.870 1.090 ;
        RECT 532.270 0.830 532.530 1.090 ;
        RECT 532.930 0.830 533.190 1.090 ;
        RECT 533.850 0.830 534.110 1.090 ;
        RECT 534.510 0.830 534.770 1.090 ;
        RECT 535.170 0.830 535.430 1.090 ;
        RECT 536.090 0.830 536.350 1.090 ;
        RECT 536.750 0.830 537.010 1.090 ;
        RECT 537.410 0.830 537.670 1.090 ;
        RECT 538.330 0.830 538.590 1.090 ;
        RECT 538.990 0.830 539.250 1.090 ;
        RECT 539.650 0.830 539.910 1.090 ;
        RECT 540.570 0.830 540.830 1.090 ;
        RECT 541.230 0.830 541.490 1.090 ;
        RECT 541.890 0.830 542.150 1.090 ;
        RECT 542.810 0.830 543.070 1.090 ;
        RECT 543.470 0.830 543.730 1.090 ;
        RECT 544.130 0.830 544.390 1.090 ;
        RECT 545.050 0.830 545.310 1.090 ;
        RECT 545.710 0.830 545.970 1.090 ;
        RECT 546.370 0.830 546.630 1.090 ;
        RECT 547.290 0.830 547.550 1.090 ;
        RECT 547.950 0.830 548.210 1.090 ;
        RECT 548.610 0.830 548.870 1.090 ;
        RECT 549.650 0.830 549.910 1.090 ;
        RECT 550.650 0.830 550.910 1.090 ;
        RECT 551.310 0.830 551.570 1.090 ;
        RECT 551.970 0.830 552.230 1.090 ;
        RECT 552.890 0.830 553.150 1.090 ;
        RECT 553.550 0.830 553.810 1.090 ;
        RECT 554.210 0.830 554.470 1.090 ;
        RECT 555.130 0.830 555.390 1.090 ;
        RECT 555.790 0.830 556.050 1.090 ;
        RECT 556.450 0.830 556.710 1.090 ;
        RECT 557.370 0.830 557.630 1.090 ;
        RECT 558.030 0.830 558.290 1.090 ;
        RECT 558.690 0.830 558.950 1.090 ;
        RECT 559.610 0.830 559.870 1.090 ;
        RECT 560.270 0.830 560.530 1.090 ;
        RECT 560.930 0.830 561.190 1.090 ;
        RECT 561.850 0.830 562.110 1.090 ;
        RECT 562.510 0.830 562.770 1.090 ;
        RECT 563.170 0.830 563.430 1.090 ;
        RECT 564.090 0.830 564.350 1.090 ;
        RECT 564.750 0.830 565.010 1.090 ;
        RECT 565.410 0.830 565.670 1.090 ;
        RECT 566.170 0.830 566.430 1.090 ;
        RECT 567.490 0.830 567.750 1.090 ;
        RECT 569.810 0.830 570.070 1.090 ;
        RECT 570.810 0.830 571.070 1.090 ;
        RECT 571.470 0.830 571.730 1.090 ;
        RECT 572.130 0.830 572.390 1.090 ;
        RECT 573.050 0.830 573.310 1.090 ;
        RECT 573.710 0.830 573.970 1.090 ;
        RECT 574.370 0.830 574.630 1.090 ;
        RECT 575.290 0.830 575.550 1.090 ;
        RECT 575.950 0.830 576.210 1.090 ;
        RECT 576.610 0.830 576.870 1.090 ;
        RECT 577.530 0.830 577.790 1.090 ;
        RECT 578.190 0.830 578.450 1.090 ;
        RECT 578.850 0.830 579.110 1.090 ;
        RECT 579.770 0.830 580.030 1.090 ;
        RECT 580.430 0.830 580.690 1.090 ;
        RECT 581.090 0.830 581.350 1.090 ;
        RECT 582.010 0.830 582.270 1.090 ;
        RECT 582.670 0.830 582.930 1.090 ;
        RECT 583.330 0.830 583.590 1.090 ;
        RECT 584.250 0.830 584.510 1.090 ;
        RECT 584.910 0.830 585.170 1.090 ;
        RECT 585.570 0.830 585.830 1.090 ;
        RECT 586.490 0.830 586.750 1.090 ;
        RECT 587.150 0.830 587.410 1.090 ;
        RECT 587.810 0.830 588.070 1.090 ;
        RECT 588.730 0.830 588.990 1.090 ;
        RECT 589.390 0.830 589.650 1.090 ;
        RECT 590.050 0.830 590.310 1.090 ;
        RECT 591.090 0.830 591.350 1.090 ;
        RECT 592.090 0.830 592.350 1.090 ;
        RECT 592.750 0.830 593.010 1.090 ;
        RECT 593.410 0.830 593.670 1.090 ;
        RECT 594.330 0.830 594.590 1.090 ;
        RECT 594.990 0.830 595.250 1.090 ;
        RECT 595.650 0.830 595.910 1.090 ;
        RECT 596.570 0.830 596.830 1.090 ;
        RECT 597.230 0.830 597.490 1.090 ;
        RECT 597.890 0.830 598.150 1.090 ;
        RECT 598.810 0.830 599.070 1.090 ;
        RECT 599.470 0.830 599.730 1.090 ;
        RECT 600.130 0.830 600.390 1.090 ;
        RECT 601.050 0.830 601.310 1.090 ;
        RECT 601.710 0.830 601.970 1.090 ;
        RECT 602.370 0.830 602.630 1.090 ;
        RECT 603.290 0.830 603.550 1.090 ;
        RECT 603.950 0.830 604.210 1.090 ;
        RECT 604.610 0.830 604.870 1.090 ;
        RECT 605.530 0.830 605.790 1.090 ;
        RECT 606.190 0.830 606.450 1.090 ;
        RECT 606.850 0.830 607.110 1.090 ;
        RECT 607.610 0.830 607.870 1.090 ;
        RECT 608.930 0.830 609.190 1.090 ;
        RECT 611.250 0.830 611.510 1.090 ;
        RECT 612.250 0.830 612.510 1.090 ;
        RECT 612.910 0.830 613.170 1.090 ;
        RECT 613.570 0.830 613.830 1.090 ;
        RECT 614.490 0.830 614.750 1.090 ;
        RECT 615.150 0.830 615.410 1.090 ;
        RECT 615.810 0.830 616.070 1.090 ;
        RECT 616.730 0.830 616.990 1.090 ;
        RECT 617.390 0.830 617.650 1.090 ;
        RECT 618.050 0.830 618.310 1.090 ;
        RECT 618.970 0.830 619.230 1.090 ;
        RECT 619.630 0.830 619.890 1.090 ;
        RECT 620.290 0.830 620.550 1.090 ;
        RECT 621.210 0.830 621.470 1.090 ;
        RECT 621.870 0.830 622.130 1.090 ;
        RECT 622.530 0.830 622.790 1.090 ;
        RECT 623.450 0.830 623.710 1.090 ;
        RECT 624.110 0.830 624.370 1.090 ;
        RECT 624.770 0.830 625.030 1.090 ;
        RECT 625.690 0.830 625.950 1.090 ;
        RECT 626.350 0.830 626.610 1.090 ;
        RECT 627.010 0.830 627.270 1.090 ;
        RECT 627.930 0.830 628.190 1.090 ;
        RECT 628.590 0.830 628.850 1.090 ;
        RECT 629.250 0.830 629.510 1.090 ;
        RECT 630.170 0.830 630.430 1.090 ;
        RECT 630.830 0.830 631.090 1.090 ;
        RECT 631.490 0.830 631.750 1.090 ;
        RECT 632.530 0.830 632.790 1.090 ;
        RECT 633.530 0.830 633.790 1.090 ;
        RECT 634.190 0.830 634.450 1.090 ;
        RECT 634.850 0.830 635.110 1.090 ;
        RECT 635.770 0.830 636.030 1.090 ;
        RECT 636.430 0.830 636.690 1.090 ;
        RECT 637.090 0.830 637.350 1.090 ;
        RECT 638.010 0.830 638.270 1.090 ;
        RECT 638.670 0.830 638.930 1.090 ;
        RECT 639.330 0.830 639.590 1.090 ;
        RECT 640.250 0.830 640.510 1.090 ;
        RECT 640.910 0.830 641.170 1.090 ;
        RECT 641.570 0.830 641.830 1.090 ;
        RECT 642.490 0.830 642.750 1.090 ;
        RECT 643.150 0.830 643.410 1.090 ;
        RECT 643.810 0.830 644.070 1.090 ;
        RECT 644.730 0.830 644.990 1.090 ;
        RECT 645.390 0.830 645.650 1.090 ;
        RECT 646.050 0.830 646.310 1.090 ;
        RECT 646.970 0.830 647.230 1.090 ;
        RECT 647.630 0.830 647.890 1.090 ;
        RECT 648.290 0.830 648.550 1.090 ;
        RECT 649.210 0.830 649.470 1.090 ;
        RECT 649.870 0.830 650.130 1.090 ;
        RECT 650.530 0.830 650.790 1.090 ;
        RECT 651.290 0.830 651.550 1.090 ;
        RECT 652.610 0.830 652.870 1.090 ;
        RECT 654.930 0.830 655.190 1.090 ;
        RECT 655.930 0.830 656.190 1.090 ;
        RECT 656.590 0.830 656.850 1.090 ;
        RECT 657.250 0.830 657.510 1.090 ;
        RECT 658.170 0.830 658.430 1.090 ;
        RECT 658.830 0.830 659.090 1.090 ;
        RECT 659.490 0.830 659.750 1.090 ;
        RECT 660.410 0.830 660.670 1.090 ;
        RECT 661.070 0.830 661.330 1.090 ;
        RECT 661.730 0.830 661.990 1.090 ;
        RECT 662.650 0.830 662.910 1.090 ;
        RECT 663.310 0.830 663.570 1.090 ;
        RECT 663.970 0.830 664.230 1.090 ;
        RECT 664.890 0.830 665.150 1.090 ;
        RECT 665.550 0.830 665.810 1.090 ;
        RECT 666.210 0.830 666.470 1.090 ;
        RECT 667.130 0.830 667.390 1.090 ;
        RECT 667.790 0.830 668.050 1.090 ;
        RECT 668.450 0.830 668.710 1.090 ;
        RECT 669.370 0.830 669.630 1.090 ;
        RECT 670.030 0.830 670.290 1.090 ;
        RECT 670.690 0.830 670.950 1.090 ;
        RECT 671.610 0.830 671.870 1.090 ;
        RECT 672.270 0.830 672.530 1.090 ;
        RECT 672.930 0.830 673.190 1.090 ;
        RECT 673.850 0.830 674.110 1.090 ;
        RECT 674.510 0.830 674.770 1.090 ;
        RECT 675.170 0.830 675.430 1.090 ;
        RECT 676.210 0.830 676.470 1.090 ;
        RECT 677.210 0.830 677.470 1.090 ;
        RECT 677.870 0.830 678.130 1.090 ;
        RECT 678.530 0.830 678.790 1.090 ;
        RECT 679.550 0.830 679.810 1.090 ;
      LAYER Metal2 ;
              RECT 3.905 11.185 8.285 17.775 ;
        RECT 14.281 11.185 18.661 17.775 ;
        RECT 24.657 11.185 29.037 17.775 ;
        RECT 35.033 11.185 39.413 17.775 ;
        RECT 46.409 11.185 50.789 17.775 ;
        RECT 56.785 11.185 61.165 17.775 ;
        RECT 67.161 11.185 71.541 17.775 ;
        RECT 77.537 11.185 81.917 17.775 ;
        RECT 88.913 11.185 93.293 17.775 ;
        RECT 99.289 11.185 103.669 17.775 ;
        RECT 109.665 11.185 114.045 17.775 ;
        RECT 120.041 11.185 124.421 17.775 ;
        RECT 131.417 11.185 135.797 17.775 ;
        RECT 141.793 11.185 146.173 17.775 ;
        RECT 152.169 11.185 156.549 17.775 ;
        RECT 162.545 11.185 166.925 17.775 ;
        RECT 173.921 11.185 178.301 17.775 ;
        RECT 184.297 11.185 188.677 17.775 ;
        RECT 194.673 11.185 199.053 17.775 ;
        RECT 205.049 11.185 209.429 17.775 ;
        RECT 216.425 11.185 220.805 17.775 ;
        RECT 226.801 11.185 231.181 17.775 ;
        RECT 237.177 11.185 241.557 17.775 ;
        RECT 247.553 11.185 251.933 17.775 ;
        RECT 258.929 11.185 263.309 17.775 ;
        RECT 269.305 11.185 273.685 17.775 ;
        RECT 279.681 11.185 284.061 17.775 ;
        RECT 290.057 11.185 294.437 17.775 ;
        RECT 301.433 11.185 305.813 17.775 ;
        RECT 311.809 11.185 316.189 17.775 ;
        RECT 322.185 11.185 326.565 17.775 ;
        RECT 332.561 11.185 336.941 17.775 ;
        RECT 343.937 11.185 348.317 17.775 ;
        RECT 354.313 11.185 358.693 17.775 ;
        RECT 364.689 11.185 369.069 17.775 ;
        RECT 375.065 11.185 379.445 17.775 ;
        RECT 386.441 11.185 390.821 17.775 ;
        RECT 396.817 11.185 401.197 17.775 ;
        RECT 407.193 11.185 411.573 17.775 ;
        RECT 417.569 11.185 421.949 17.775 ;
        RECT 428.945 11.185 433.325 17.775 ;
        RECT 439.321 11.185 443.701 17.775 ;
        RECT 449.697 11.185 454.077 17.775 ;
        RECT 460.073 11.185 464.453 17.775 ;
        RECT 471.449 11.185 475.829 17.775 ;
        RECT 481.825 11.185 486.205 17.775 ;
        RECT 492.201 11.185 496.581 17.775 ;
        RECT 502.577 11.185 506.957 17.775 ;
        RECT 513.953 11.185 518.333 17.775 ;
        RECT 524.329 11.185 528.709 17.775 ;
        RECT 534.705 11.185 539.085 17.775 ;
        RECT 545.081 11.185 549.461 17.775 ;
        RECT 556.457 11.185 560.837 17.775 ;
        RECT 566.833 11.185 571.213 17.775 ;
        RECT 577.209 11.185 581.589 17.775 ;
        RECT 587.585 11.185 591.965 17.775 ;
        RECT 598.961 11.185 603.341 17.775 ;
        RECT 609.337 11.185 613.717 17.775 ;
        RECT 619.713 11.185 624.093 17.775 ;
        RECT 630.089 11.185 634.469 17.775 ;
        RECT 641.465 11.185 645.845 17.775 ;
        RECT 651.841 11.185 656.221 17.775 ;
        RECT 662.217 11.185 666.597 17.775 ;
        RECT 672.593 11.185 676.973 17.775 ;
        RECT 3.915 49.781 8.295 56.371 ;
        RECT 14.291 49.781 18.671 56.371 ;
        RECT 24.667 49.781 29.047 56.371 ;
        RECT 35.043 49.781 39.423 56.371 ;
        RECT 46.419 49.781 50.799 56.371 ;
        RECT 56.795 49.781 61.175 56.371 ;
        RECT 67.171 49.781 71.551 56.371 ;
        RECT 77.547 49.781 81.927 56.371 ;
        RECT 88.923 49.781 93.303 56.371 ;
        RECT 99.299 49.781 103.679 56.371 ;
        RECT 109.675 49.781 114.055 56.371 ;
        RECT 120.051 49.781 124.431 56.371 ;
        RECT 131.427 49.781 135.807 56.371 ;
        RECT 141.803 49.781 146.183 56.371 ;
        RECT 152.179 49.781 156.559 56.371 ;
        RECT 162.555 49.781 166.935 56.371 ;
        RECT 173.931 49.781 178.311 56.371 ;
        RECT 184.307 49.781 188.687 56.371 ;
        RECT 194.683 49.781 199.063 56.371 ;
        RECT 205.059 49.781 209.439 56.371 ;
        RECT 216.435 49.781 220.815 56.371 ;
        RECT 226.811 49.781 231.191 56.371 ;
        RECT 237.187 49.781 241.567 56.371 ;
        RECT 247.563 49.781 251.943 56.371 ;
        RECT 258.939 49.781 263.319 56.371 ;
        RECT 269.315 49.781 273.695 56.371 ;
        RECT 279.691 49.781 284.071 56.371 ;
        RECT 290.067 49.781 294.447 56.371 ;
        RECT 301.443 49.781 305.823 56.371 ;
        RECT 311.819 49.781 316.199 56.371 ;
        RECT 322.195 49.781 326.575 56.371 ;
        RECT 332.571 49.781 336.951 56.371 ;
        RECT 343.947 49.781 348.327 56.371 ;
        RECT 354.323 49.781 358.703 56.371 ;
        RECT 364.699 49.781 369.079 56.371 ;
        RECT 375.075 49.781 379.455 56.371 ;
        RECT 386.451 49.781 390.831 56.371 ;
        RECT 396.827 49.781 401.207 56.371 ;
        RECT 407.203 49.781 411.583 56.371 ;
        RECT 417.579 49.781 421.959 56.371 ;
        RECT 428.955 49.781 433.335 56.371 ;
        RECT 439.331 49.781 443.711 56.371 ;
        RECT 449.707 49.781 454.087 56.371 ;
        RECT 460.083 49.781 464.463 56.371 ;
        RECT 471.459 49.781 475.839 56.371 ;
        RECT 481.835 49.781 486.215 56.371 ;
        RECT 492.211 49.781 496.591 56.371 ;
        RECT 502.587 49.781 506.967 56.371 ;
        RECT 513.963 49.781 518.343 56.371 ;
        RECT 524.339 49.781 528.719 56.371 ;
        RECT 534.715 49.781 539.095 56.371 ;
        RECT 545.091 49.781 549.471 56.371 ;
        RECT 556.467 49.781 560.847 56.371 ;
        RECT 566.843 49.781 571.223 56.371 ;
        RECT 577.219 49.781 581.599 56.371 ;
        RECT 587.595 49.781 591.975 56.371 ;
        RECT 598.971 49.781 603.351 56.371 ;
        RECT 609.347 49.781 613.727 56.371 ;
        RECT 619.723 49.781 624.103 56.371 ;
        RECT 630.099 49.781 634.479 56.371 ;
        RECT 641.475 49.781 645.855 56.371 ;
        RECT 651.851 49.781 656.231 56.371 ;
        RECT 662.227 49.781 666.607 56.371 ;
        RECT 672.603 49.781 676.983 56.371 ;

        RECT 1.975 59.890 41.085 60.305 ;
        RECT 44.545 59.890 83.655 60.305 ;
        RECT 87.115 59.890 126.225 60.305 ;
        RECT 129.685 59.890 168.795 60.305 ;
        RECT 172.255 59.890 211.365 60.305 ;
        RECT 214.825 59.890 253.935 60.305 ;
        RECT 257.395 59.890 296.505 60.305 ;
        RECT 299.965 59.890 339.075 60.305 ;
        RECT 342.535 59.890 381.645 60.305 ;
        RECT 385.105 59.890 424.215 60.305 ;
        RECT 427.675 59.890 466.785 60.305 ;
        RECT 470.245 59.890 509.355 60.305 ;
        RECT 512.815 59.890 551.925 60.305 ;
        RECT 555.385 59.890 594.495 60.305 ;
        RECT 597.955 59.890 637.065 60.305 ;
        RECT 640.525 59.890 679.635 60.305 ;
        RECT 0.765 58.745 1.145 59.125 ;
        RECT 0.765 58.085 1.145 58.465 ;
        RECT 0.765 57.425 1.145 57.805 ;
        RECT 0.765 56.765 1.145 57.145 ;
        RECT 0.765 56.105 1.145 56.485 ;
        RECT 0.765 55.445 1.145 55.825 ;
        RECT 0.765 54.785 1.145 55.165 ;
        RECT 0.765 54.125 1.145 54.505 ;
        RECT 0.765 53.465 1.145 53.845 ;
        RECT 0.765 52.805 1.145 53.185 ;
        RECT 0.765 52.145 1.145 52.525 ;
        RECT 0.765 51.485 1.145 51.865 ;
        RECT 0.765 50.825 1.145 51.205 ;
        RECT 0.765 50.165 1.145 50.545 ;
        RECT 5.250 47.805 5.630 48.185 ;
        RECT 5.910 47.805 6.290 48.185 ;
        RECT 6.570 47.805 6.950 48.185 ;
        RECT 5.250 47.145 5.630 47.525 ;
        RECT 5.910 47.145 6.290 47.525 ;
        RECT 6.570 47.145 6.950 47.525 ;
        RECT 5.250 46.485 5.630 46.865 ;
        RECT 5.910 46.485 6.290 46.865 ;
        RECT 6.570 46.485 6.950 46.865 ;
        RECT 5.250 22.205 5.630 22.585 ;
        RECT 5.910 22.205 6.290 22.585 ;
        RECT 6.570 22.205 6.950 22.585 ;
        RECT 5.250 21.545 5.630 21.925 ;
        RECT 5.910 21.545 6.290 21.925 ;
        RECT 6.570 21.545 6.950 21.925 ;
        RECT 5.250 20.885 5.630 21.265 ;
        RECT 5.910 20.885 6.290 21.265 ;
        RECT 6.570 20.885 6.950 21.265 ;
        RECT 9.000 9.150 9.525 59.890 ;
        RECT 11.055 58.745 11.435 59.125 ;
        RECT 11.055 58.085 11.435 58.465 ;
        RECT 11.055 57.425 11.435 57.805 ;
        RECT 11.055 56.765 11.435 57.145 ;
        RECT 11.055 56.105 11.435 56.485 ;
        RECT 11.055 55.445 11.435 55.825 ;
        RECT 11.055 54.785 11.435 55.165 ;
        RECT 11.055 54.125 11.435 54.505 ;
        RECT 11.055 53.465 11.435 53.845 ;
        RECT 11.055 52.805 11.435 53.185 ;
        RECT 11.055 52.145 11.435 52.525 ;
        RECT 11.055 51.485 11.435 51.865 ;
        RECT 11.055 50.825 11.435 51.205 ;
        RECT 11.055 50.165 11.435 50.545 ;
        RECT 12.440 9.150 12.965 59.890 ;
        RECT 21.340 58.745 21.720 59.125 ;
        RECT 21.340 58.085 21.720 58.465 ;
        RECT 21.340 57.425 21.720 57.805 ;
        RECT 21.340 56.765 21.720 57.145 ;
        RECT 21.340 56.105 21.720 56.485 ;
        RECT 21.340 55.445 21.720 55.825 ;
        RECT 21.340 54.785 21.720 55.165 ;
        RECT 21.340 54.125 21.720 54.505 ;
        RECT 21.340 53.465 21.720 53.845 ;
        RECT 21.340 52.805 21.720 53.185 ;
        RECT 21.340 52.145 21.720 52.525 ;
        RECT 21.340 51.485 21.720 51.865 ;
        RECT 21.340 50.825 21.720 51.205 ;
        RECT 21.340 50.165 21.720 50.545 ;
        RECT 15.550 45.105 15.930 45.485 ;
        RECT 16.210 45.105 16.590 45.485 ;
        RECT 16.870 45.105 17.250 45.485 ;
        RECT 15.550 44.445 15.930 44.825 ;
        RECT 16.210 44.445 16.590 44.825 ;
        RECT 16.870 44.445 17.250 44.825 ;
        RECT 15.550 43.785 15.930 44.165 ;
        RECT 16.210 43.785 16.590 44.165 ;
        RECT 16.870 43.785 17.250 44.165 ;
        RECT 25.825 42.405 26.205 42.785 ;
        RECT 26.485 42.405 26.865 42.785 ;
        RECT 27.145 42.405 27.525 42.785 ;
        RECT 25.825 41.745 26.205 42.125 ;
        RECT 26.485 41.745 26.865 42.125 ;
        RECT 27.145 41.745 27.525 42.125 ;
        RECT 25.825 41.085 26.205 41.465 ;
        RECT 26.485 41.085 26.865 41.465 ;
        RECT 27.145 41.085 27.525 41.465 ;
        RECT 25.825 27.605 26.205 27.985 ;
        RECT 26.485 27.605 26.865 27.985 ;
        RECT 27.145 27.605 27.525 27.985 ;
        RECT 25.825 26.945 26.205 27.325 ;
        RECT 26.485 26.945 26.865 27.325 ;
        RECT 27.145 26.945 27.525 27.325 ;
        RECT 25.825 26.285 26.205 26.665 ;
        RECT 26.485 26.285 26.865 26.665 ;
        RECT 27.145 26.285 27.525 26.665 ;
        RECT 15.550 24.905 15.930 25.285 ;
        RECT 16.210 24.905 16.590 25.285 ;
        RECT 16.870 24.905 17.250 25.285 ;
        RECT 15.550 24.245 15.930 24.625 ;
        RECT 16.210 24.245 16.590 24.625 ;
        RECT 16.870 24.245 17.250 24.625 ;
        RECT 15.550 23.585 15.930 23.965 ;
        RECT 16.210 23.585 16.590 23.965 ;
        RECT 16.870 23.585 17.250 23.965 ;
        RECT 9.000 9.100 12.965 9.150 ;
        RECT 29.575 9.150 30.100 59.890 ;
        RECT 31.630 58.745 32.010 59.125 ;
        RECT 31.630 58.085 32.010 58.465 ;
        RECT 31.630 57.425 32.010 57.805 ;
        RECT 31.630 56.765 32.010 57.145 ;
        RECT 31.630 56.105 32.010 56.485 ;
        RECT 31.630 55.445 32.010 55.825 ;
        RECT 31.630 54.785 32.010 55.165 ;
        RECT 31.630 54.125 32.010 54.505 ;
        RECT 31.630 53.465 32.010 53.845 ;
        RECT 31.630 52.805 32.010 53.185 ;
        RECT 31.630 52.145 32.010 52.525 ;
        RECT 31.630 51.485 32.010 51.865 ;
        RECT 31.630 50.825 32.010 51.205 ;
        RECT 31.630 50.165 32.010 50.545 ;
        RECT 33.015 9.150 33.540 59.890 ;
        RECT 41.915 58.745 42.295 59.125 ;
        RECT 43.335 58.745 43.715 59.125 ;
        RECT 41.915 58.085 42.295 58.465 ;
        RECT 43.335 58.085 43.715 58.465 ;
        RECT 41.915 57.425 42.295 57.805 ;
        RECT 43.335 57.425 43.715 57.805 ;
        RECT 41.915 56.765 42.295 57.145 ;
        RECT 43.335 56.765 43.715 57.145 ;
        RECT 41.915 56.105 42.295 56.485 ;
        RECT 43.335 56.105 43.715 56.485 ;
        RECT 41.915 55.445 42.295 55.825 ;
        RECT 43.335 55.445 43.715 55.825 ;
        RECT 41.915 54.785 42.295 55.165 ;
        RECT 43.335 54.785 43.715 55.165 ;
        RECT 41.915 54.125 42.295 54.505 ;
        RECT 43.335 54.125 43.715 54.505 ;
        RECT 41.915 53.465 42.295 53.845 ;
        RECT 43.335 53.465 43.715 53.845 ;
        RECT 41.915 52.805 42.295 53.185 ;
        RECT 43.335 52.805 43.715 53.185 ;
        RECT 41.915 52.145 42.295 52.525 ;
        RECT 43.335 52.145 43.715 52.525 ;
        RECT 41.915 51.485 42.295 51.865 ;
        RECT 43.335 51.485 43.715 51.865 ;
        RECT 41.915 50.825 42.295 51.205 ;
        RECT 43.335 50.825 43.715 51.205 ;
        RECT 41.915 50.165 42.295 50.545 ;
        RECT 43.335 50.165 43.715 50.545 ;
        RECT 47.820 47.805 48.200 48.185 ;
        RECT 48.480 47.805 48.860 48.185 ;
        RECT 49.140 47.805 49.520 48.185 ;
        RECT 47.820 47.145 48.200 47.525 ;
        RECT 48.480 47.145 48.860 47.525 ;
        RECT 49.140 47.145 49.520 47.525 ;
        RECT 47.820 46.485 48.200 46.865 ;
        RECT 48.480 46.485 48.860 46.865 ;
        RECT 49.140 46.485 49.520 46.865 ;
        RECT 36.125 39.705 36.505 40.085 ;
        RECT 36.785 39.705 37.165 40.085 ;
        RECT 37.445 39.705 37.825 40.085 ;
        RECT 36.125 39.045 36.505 39.425 ;
        RECT 36.785 39.045 37.165 39.425 ;
        RECT 37.445 39.045 37.825 39.425 ;
        RECT 36.125 38.385 36.505 38.765 ;
        RECT 36.785 38.385 37.165 38.765 ;
        RECT 37.445 38.385 37.825 38.765 ;
        RECT 36.125 30.305 36.505 30.685 ;
        RECT 36.785 30.305 37.165 30.685 ;
        RECT 37.445 30.305 37.825 30.685 ;
        RECT 36.125 29.645 36.505 30.025 ;
        RECT 36.785 29.645 37.165 30.025 ;
        RECT 37.445 29.645 37.825 30.025 ;
        RECT 36.125 28.985 36.505 29.365 ;
        RECT 36.785 28.985 37.165 29.365 ;
        RECT 37.445 28.985 37.825 29.365 ;
        RECT 47.820 22.205 48.200 22.585 ;
        RECT 48.480 22.205 48.860 22.585 ;
        RECT 49.140 22.205 49.520 22.585 ;
        RECT 47.820 21.545 48.200 21.925 ;
        RECT 48.480 21.545 48.860 21.925 ;
        RECT 49.140 21.545 49.520 21.925 ;
        RECT 47.820 20.885 48.200 21.265 ;
        RECT 48.480 20.885 48.860 21.265 ;
        RECT 49.140 20.885 49.520 21.265 ;
        RECT 9.000 8.770 20.385 9.100 ;
        RECT 9.000 8.750 12.965 8.770 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 0.850 4.690 1.230 5.070 ;
        RECT 1.990 4.690 2.370 5.070 ;
        RECT 8.030 4.720 8.410 5.100 ;
        RECT 8.690 4.720 9.070 5.100 ;
        RECT 9.350 4.720 9.730 5.100 ;
        RECT 14.560 4.690 14.940 5.070 ;
        RECT 15.220 4.690 15.600 5.070 ;
        RECT 15.880 4.690 16.260 5.070 ;
        RECT 17.920 4.690 18.300 5.070 ;
        RECT 18.580 4.690 18.960 5.070 ;
        RECT 19.240 4.690 19.620 5.070 ;
        RECT 3.490 2.950 3.860 4.550 ;
        RECT 20.055 4.150 20.385 8.770 ;
        RECT 29.575 8.750 33.540 9.150 ;
        RECT 51.570 9.150 52.095 59.890 ;
        RECT 53.625 58.745 54.005 59.125 ;
        RECT 53.625 58.085 54.005 58.465 ;
        RECT 53.625 57.425 54.005 57.805 ;
        RECT 53.625 56.765 54.005 57.145 ;
        RECT 53.625 56.105 54.005 56.485 ;
        RECT 53.625 55.445 54.005 55.825 ;
        RECT 53.625 54.785 54.005 55.165 ;
        RECT 53.625 54.125 54.005 54.505 ;
        RECT 53.625 53.465 54.005 53.845 ;
        RECT 53.625 52.805 54.005 53.185 ;
        RECT 53.625 52.145 54.005 52.525 ;
        RECT 53.625 51.485 54.005 51.865 ;
        RECT 53.625 50.825 54.005 51.205 ;
        RECT 53.625 50.165 54.005 50.545 ;
        RECT 55.010 9.150 55.535 59.890 ;
        RECT 63.910 58.745 64.290 59.125 ;
        RECT 63.910 58.085 64.290 58.465 ;
        RECT 63.910 57.425 64.290 57.805 ;
        RECT 63.910 56.765 64.290 57.145 ;
        RECT 63.910 56.105 64.290 56.485 ;
        RECT 63.910 55.445 64.290 55.825 ;
        RECT 63.910 54.785 64.290 55.165 ;
        RECT 63.910 54.125 64.290 54.505 ;
        RECT 63.910 53.465 64.290 53.845 ;
        RECT 63.910 52.805 64.290 53.185 ;
        RECT 63.910 52.145 64.290 52.525 ;
        RECT 63.910 51.485 64.290 51.865 ;
        RECT 63.910 50.825 64.290 51.205 ;
        RECT 63.910 50.165 64.290 50.545 ;
        RECT 58.120 45.105 58.500 45.485 ;
        RECT 58.780 45.105 59.160 45.485 ;
        RECT 59.440 45.105 59.820 45.485 ;
        RECT 58.120 44.445 58.500 44.825 ;
        RECT 58.780 44.445 59.160 44.825 ;
        RECT 59.440 44.445 59.820 44.825 ;
        RECT 58.120 43.785 58.500 44.165 ;
        RECT 58.780 43.785 59.160 44.165 ;
        RECT 59.440 43.785 59.820 44.165 ;
        RECT 68.395 42.405 68.775 42.785 ;
        RECT 69.055 42.405 69.435 42.785 ;
        RECT 69.715 42.405 70.095 42.785 ;
        RECT 68.395 41.745 68.775 42.125 ;
        RECT 69.055 41.745 69.435 42.125 ;
        RECT 69.715 41.745 70.095 42.125 ;
        RECT 68.395 41.085 68.775 41.465 ;
        RECT 69.055 41.085 69.435 41.465 ;
        RECT 69.715 41.085 70.095 41.465 ;
        RECT 68.395 27.605 68.775 27.985 ;
        RECT 69.055 27.605 69.435 27.985 ;
        RECT 69.715 27.605 70.095 27.985 ;
        RECT 68.395 26.945 68.775 27.325 ;
        RECT 69.055 26.945 69.435 27.325 ;
        RECT 69.715 26.945 70.095 27.325 ;
        RECT 68.395 26.285 68.775 26.665 ;
        RECT 69.055 26.285 69.435 26.665 ;
        RECT 69.715 26.285 70.095 26.665 ;
        RECT 58.120 24.905 58.500 25.285 ;
        RECT 58.780 24.905 59.160 25.285 ;
        RECT 59.440 24.905 59.820 25.285 ;
        RECT 58.120 24.245 58.500 24.625 ;
        RECT 58.780 24.245 59.160 24.625 ;
        RECT 59.440 24.245 59.820 24.625 ;
        RECT 58.120 23.585 58.500 23.965 ;
        RECT 58.780 23.585 59.160 23.965 ;
        RECT 59.440 23.585 59.820 23.965 ;
        RECT 51.570 9.100 55.535 9.150 ;
        RECT 72.145 9.150 72.670 59.890 ;
        RECT 74.200 58.745 74.580 59.125 ;
        RECT 74.200 58.085 74.580 58.465 ;
        RECT 74.200 57.425 74.580 57.805 ;
        RECT 74.200 56.765 74.580 57.145 ;
        RECT 74.200 56.105 74.580 56.485 ;
        RECT 74.200 55.445 74.580 55.825 ;
        RECT 74.200 54.785 74.580 55.165 ;
        RECT 74.200 54.125 74.580 54.505 ;
        RECT 74.200 53.465 74.580 53.845 ;
        RECT 74.200 52.805 74.580 53.185 ;
        RECT 74.200 52.145 74.580 52.525 ;
        RECT 74.200 51.485 74.580 51.865 ;
        RECT 74.200 50.825 74.580 51.205 ;
        RECT 74.200 50.165 74.580 50.545 ;
        RECT 75.585 9.150 76.110 59.890 ;
        RECT 84.485 58.745 84.865 59.125 ;
        RECT 85.905 58.745 86.285 59.125 ;
        RECT 84.485 58.085 84.865 58.465 ;
        RECT 85.905 58.085 86.285 58.465 ;
        RECT 84.485 57.425 84.865 57.805 ;
        RECT 85.905 57.425 86.285 57.805 ;
        RECT 84.485 56.765 84.865 57.145 ;
        RECT 85.905 56.765 86.285 57.145 ;
        RECT 84.485 56.105 84.865 56.485 ;
        RECT 85.905 56.105 86.285 56.485 ;
        RECT 84.485 55.445 84.865 55.825 ;
        RECT 85.905 55.445 86.285 55.825 ;
        RECT 84.485 54.785 84.865 55.165 ;
        RECT 85.905 54.785 86.285 55.165 ;
        RECT 84.485 54.125 84.865 54.505 ;
        RECT 85.905 54.125 86.285 54.505 ;
        RECT 84.485 53.465 84.865 53.845 ;
        RECT 85.905 53.465 86.285 53.845 ;
        RECT 84.485 52.805 84.865 53.185 ;
        RECT 85.905 52.805 86.285 53.185 ;
        RECT 84.485 52.145 84.865 52.525 ;
        RECT 85.905 52.145 86.285 52.525 ;
        RECT 84.485 51.485 84.865 51.865 ;
        RECT 85.905 51.485 86.285 51.865 ;
        RECT 84.485 50.825 84.865 51.205 ;
        RECT 85.905 50.825 86.285 51.205 ;
        RECT 84.485 50.165 84.865 50.545 ;
        RECT 85.905 50.165 86.285 50.545 ;
        RECT 90.390 47.805 90.770 48.185 ;
        RECT 91.050 47.805 91.430 48.185 ;
        RECT 91.710 47.805 92.090 48.185 ;
        RECT 90.390 47.145 90.770 47.525 ;
        RECT 91.050 47.145 91.430 47.525 ;
        RECT 91.710 47.145 92.090 47.525 ;
        RECT 90.390 46.485 90.770 46.865 ;
        RECT 91.050 46.485 91.430 46.865 ;
        RECT 91.710 46.485 92.090 46.865 ;
        RECT 78.695 39.705 79.075 40.085 ;
        RECT 79.355 39.705 79.735 40.085 ;
        RECT 80.015 39.705 80.395 40.085 ;
        RECT 78.695 39.045 79.075 39.425 ;
        RECT 79.355 39.045 79.735 39.425 ;
        RECT 80.015 39.045 80.395 39.425 ;
        RECT 78.695 38.385 79.075 38.765 ;
        RECT 79.355 38.385 79.735 38.765 ;
        RECT 80.015 38.385 80.395 38.765 ;
        RECT 78.695 30.305 79.075 30.685 ;
        RECT 79.355 30.305 79.735 30.685 ;
        RECT 80.015 30.305 80.395 30.685 ;
        RECT 78.695 29.645 79.075 30.025 ;
        RECT 79.355 29.645 79.735 30.025 ;
        RECT 80.015 29.645 80.395 30.025 ;
        RECT 78.695 28.985 79.075 29.365 ;
        RECT 79.355 28.985 79.735 29.365 ;
        RECT 80.015 28.985 80.395 29.365 ;
        RECT 90.390 22.205 90.770 22.585 ;
        RECT 91.050 22.205 91.430 22.585 ;
        RECT 91.710 22.205 92.090 22.585 ;
        RECT 90.390 21.545 90.770 21.925 ;
        RECT 91.050 21.545 91.430 21.925 ;
        RECT 91.710 21.545 92.090 21.925 ;
        RECT 90.390 20.885 90.770 21.265 ;
        RECT 91.050 20.885 91.430 21.265 ;
        RECT 91.710 20.885 92.090 21.265 ;
        RECT 51.570 8.770 69.355 9.100 ;
        RECT 51.570 8.750 55.535 8.770 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 38.750 8.090 39.130 8.470 ;
        RECT 53.580 8.090 53.960 8.470 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 38.750 7.430 39.130 7.810 ;
        RECT 53.580 7.430 53.960 7.810 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 38.750 6.770 39.130 7.150 ;
        RECT 53.580 6.770 53.960 7.150 ;
        RECT 26.220 4.720 26.600 5.100 ;
        RECT 26.880 4.720 27.260 5.100 ;
        RECT 27.540 4.720 27.920 5.100 ;
        RECT 32.750 4.690 33.130 5.070 ;
        RECT 33.410 4.690 33.790 5.070 ;
        RECT 34.070 4.690 34.450 5.070 ;
        RECT 36.130 4.690 36.510 5.070 ;
        RECT 42.170 4.720 42.550 5.100 ;
        RECT 42.830 4.720 43.210 5.100 ;
        RECT 43.490 4.720 43.870 5.100 ;
        RECT 48.700 4.690 49.080 5.070 ;
        RECT 49.360 4.690 49.740 5.070 ;
        RECT 50.020 4.690 50.400 5.070 ;
        RECT 57.000 4.720 57.380 5.100 ;
        RECT 57.660 4.720 58.040 5.100 ;
        RECT 58.320 4.720 58.700 5.100 ;
        RECT 63.530 4.690 63.910 5.070 ;
        RECT 64.190 4.690 64.570 5.070 ;
        RECT 64.850 4.690 65.230 5.070 ;
        RECT 66.890 4.690 67.270 5.070 ;
        RECT 67.550 4.690 67.930 5.070 ;
        RECT 68.210 4.690 68.590 5.070 ;
        RECT 4.170 3.420 4.550 3.800 ;
        RECT 20.030 3.770 20.410 4.150 ;
        RECT 3.490 2.580 4.190 2.950 ;
        RECT 4.580 2.760 4.960 3.140 ;
        RECT 6.995 2.950 10.205 3.300 ;
        RECT 3.820 2.305 4.190 2.580 ;
        RECT 6.995 2.305 7.345 2.950 ;
        RECT 11.480 2.760 13.000 3.255 ;
        RECT 14.945 3.125 15.325 3.150 ;
        RECT 13.865 2.795 15.325 3.125 ;
        RECT 11.480 2.600 11.890 2.760 ;
        RECT 3.820 1.955 7.345 2.305 ;
        RECT 7.645 2.250 11.890 2.600 ;
        RECT 12.090 1.885 12.470 1.910 ;
        RECT 13.865 1.885 14.195 2.795 ;
        RECT 14.945 2.770 15.325 2.795 ;
        RECT 21.680 2.950 22.050 4.550 ;
        RECT 22.360 3.420 22.740 3.800 ;
        RECT 21.680 2.580 22.380 2.950 ;
        RECT 22.770 2.760 23.150 3.140 ;
        RECT 25.185 2.950 28.395 3.300 ;
        RECT 22.010 2.305 22.380 2.580 ;
        RECT 25.185 2.305 25.535 2.950 ;
        RECT 29.670 2.760 31.190 3.255 ;
        RECT 33.135 3.125 33.515 3.150 ;
        RECT 32.055 2.795 33.515 3.125 ;
        RECT 29.670 2.600 30.080 2.760 ;
        RECT 22.010 1.955 25.535 2.305 ;
        RECT 25.835 2.250 30.080 2.600 ;
        RECT 12.090 1.555 14.195 1.885 ;
        RECT 30.280 1.885 30.660 1.910 ;
        RECT 32.055 1.885 32.385 2.795 ;
        RECT 33.135 2.770 33.515 2.795 ;
        RECT 37.630 2.950 38.000 4.550 ;
        RECT 38.310 3.420 38.690 3.800 ;
        RECT 37.630 2.580 38.330 2.950 ;
        RECT 38.720 2.760 39.100 3.140 ;
        RECT 41.135 2.950 44.345 3.300 ;
        RECT 37.960 2.305 38.330 2.580 ;
        RECT 41.135 2.305 41.485 2.950 ;
        RECT 45.620 2.760 47.140 3.255 ;
        RECT 49.085 3.125 49.465 3.150 ;
        RECT 48.005 2.795 49.465 3.125 ;
        RECT 45.620 2.600 46.030 2.760 ;
        RECT 37.960 1.955 41.485 2.305 ;
        RECT 41.785 2.250 46.030 2.600 ;
        RECT 30.280 1.555 32.385 1.885 ;
        RECT 46.230 1.885 46.610 1.910 ;
        RECT 48.005 1.885 48.335 2.795 ;
        RECT 49.085 2.770 49.465 2.795 ;
        RECT 52.460 2.950 52.830 4.550 ;
        RECT 69.025 4.150 69.355 8.770 ;
        RECT 72.145 8.750 76.110 9.150 ;
        RECT 94.140 9.150 94.665 59.890 ;
        RECT 96.195 58.745 96.575 59.125 ;
        RECT 96.195 58.085 96.575 58.465 ;
        RECT 96.195 57.425 96.575 57.805 ;
        RECT 96.195 56.765 96.575 57.145 ;
        RECT 96.195 56.105 96.575 56.485 ;
        RECT 96.195 55.445 96.575 55.825 ;
        RECT 96.195 54.785 96.575 55.165 ;
        RECT 96.195 54.125 96.575 54.505 ;
        RECT 96.195 53.465 96.575 53.845 ;
        RECT 96.195 52.805 96.575 53.185 ;
        RECT 96.195 52.145 96.575 52.525 ;
        RECT 96.195 51.485 96.575 51.865 ;
        RECT 96.195 50.825 96.575 51.205 ;
        RECT 96.195 50.165 96.575 50.545 ;
        RECT 97.580 9.150 98.105 59.890 ;
        RECT 106.480 58.745 106.860 59.125 ;
        RECT 106.480 58.085 106.860 58.465 ;
        RECT 106.480 57.425 106.860 57.805 ;
        RECT 106.480 56.765 106.860 57.145 ;
        RECT 106.480 56.105 106.860 56.485 ;
        RECT 106.480 55.445 106.860 55.825 ;
        RECT 106.480 54.785 106.860 55.165 ;
        RECT 106.480 54.125 106.860 54.505 ;
        RECT 106.480 53.465 106.860 53.845 ;
        RECT 106.480 52.805 106.860 53.185 ;
        RECT 106.480 52.145 106.860 52.525 ;
        RECT 106.480 51.485 106.860 51.865 ;
        RECT 106.480 50.825 106.860 51.205 ;
        RECT 106.480 50.165 106.860 50.545 ;
        RECT 100.690 45.105 101.070 45.485 ;
        RECT 101.350 45.105 101.730 45.485 ;
        RECT 102.010 45.105 102.390 45.485 ;
        RECT 100.690 44.445 101.070 44.825 ;
        RECT 101.350 44.445 101.730 44.825 ;
        RECT 102.010 44.445 102.390 44.825 ;
        RECT 100.690 43.785 101.070 44.165 ;
        RECT 101.350 43.785 101.730 44.165 ;
        RECT 102.010 43.785 102.390 44.165 ;
        RECT 110.965 42.405 111.345 42.785 ;
        RECT 111.625 42.405 112.005 42.785 ;
        RECT 112.285 42.405 112.665 42.785 ;
        RECT 110.965 41.745 111.345 42.125 ;
        RECT 111.625 41.745 112.005 42.125 ;
        RECT 112.285 41.745 112.665 42.125 ;
        RECT 110.965 41.085 111.345 41.465 ;
        RECT 111.625 41.085 112.005 41.465 ;
        RECT 112.285 41.085 112.665 41.465 ;
        RECT 110.965 27.605 111.345 27.985 ;
        RECT 111.625 27.605 112.005 27.985 ;
        RECT 112.285 27.605 112.665 27.985 ;
        RECT 110.965 26.945 111.345 27.325 ;
        RECT 111.625 26.945 112.005 27.325 ;
        RECT 112.285 26.945 112.665 27.325 ;
        RECT 110.965 26.285 111.345 26.665 ;
        RECT 111.625 26.285 112.005 26.665 ;
        RECT 112.285 26.285 112.665 26.665 ;
        RECT 100.690 24.905 101.070 25.285 ;
        RECT 101.350 24.905 101.730 25.285 ;
        RECT 102.010 24.905 102.390 25.285 ;
        RECT 100.690 24.245 101.070 24.625 ;
        RECT 101.350 24.245 101.730 24.625 ;
        RECT 102.010 24.245 102.390 24.625 ;
        RECT 100.690 23.585 101.070 23.965 ;
        RECT 101.350 23.585 101.730 23.965 ;
        RECT 102.010 23.585 102.390 23.965 ;
        RECT 94.140 9.100 98.105 9.150 ;
        RECT 114.715 9.150 115.240 59.890 ;
        RECT 116.770 58.745 117.150 59.125 ;
        RECT 116.770 58.085 117.150 58.465 ;
        RECT 116.770 57.425 117.150 57.805 ;
        RECT 116.770 56.765 117.150 57.145 ;
        RECT 116.770 56.105 117.150 56.485 ;
        RECT 116.770 55.445 117.150 55.825 ;
        RECT 116.770 54.785 117.150 55.165 ;
        RECT 116.770 54.125 117.150 54.505 ;
        RECT 116.770 53.465 117.150 53.845 ;
        RECT 116.770 52.805 117.150 53.185 ;
        RECT 116.770 52.145 117.150 52.525 ;
        RECT 116.770 51.485 117.150 51.865 ;
        RECT 116.770 50.825 117.150 51.205 ;
        RECT 116.770 50.165 117.150 50.545 ;
        RECT 118.155 9.150 118.680 59.890 ;
        RECT 127.055 58.745 127.435 59.125 ;
        RECT 128.475 58.745 128.855 59.125 ;
        RECT 127.055 58.085 127.435 58.465 ;
        RECT 128.475 58.085 128.855 58.465 ;
        RECT 127.055 57.425 127.435 57.805 ;
        RECT 128.475 57.425 128.855 57.805 ;
        RECT 127.055 56.765 127.435 57.145 ;
        RECT 128.475 56.765 128.855 57.145 ;
        RECT 127.055 56.105 127.435 56.485 ;
        RECT 128.475 56.105 128.855 56.485 ;
        RECT 127.055 55.445 127.435 55.825 ;
        RECT 128.475 55.445 128.855 55.825 ;
        RECT 127.055 54.785 127.435 55.165 ;
        RECT 128.475 54.785 128.855 55.165 ;
        RECT 127.055 54.125 127.435 54.505 ;
        RECT 128.475 54.125 128.855 54.505 ;
        RECT 127.055 53.465 127.435 53.845 ;
        RECT 128.475 53.465 128.855 53.845 ;
        RECT 127.055 52.805 127.435 53.185 ;
        RECT 128.475 52.805 128.855 53.185 ;
        RECT 127.055 52.145 127.435 52.525 ;
        RECT 128.475 52.145 128.855 52.525 ;
        RECT 127.055 51.485 127.435 51.865 ;
        RECT 128.475 51.485 128.855 51.865 ;
        RECT 127.055 50.825 127.435 51.205 ;
        RECT 128.475 50.825 128.855 51.205 ;
        RECT 127.055 50.165 127.435 50.545 ;
        RECT 128.475 50.165 128.855 50.545 ;
        RECT 132.960 47.805 133.340 48.185 ;
        RECT 133.620 47.805 134.000 48.185 ;
        RECT 134.280 47.805 134.660 48.185 ;
        RECT 132.960 47.145 133.340 47.525 ;
        RECT 133.620 47.145 134.000 47.525 ;
        RECT 134.280 47.145 134.660 47.525 ;
        RECT 132.960 46.485 133.340 46.865 ;
        RECT 133.620 46.485 134.000 46.865 ;
        RECT 134.280 46.485 134.660 46.865 ;
        RECT 121.265 39.705 121.645 40.085 ;
        RECT 121.925 39.705 122.305 40.085 ;
        RECT 122.585 39.705 122.965 40.085 ;
        RECT 121.265 39.045 121.645 39.425 ;
        RECT 121.925 39.045 122.305 39.425 ;
        RECT 122.585 39.045 122.965 39.425 ;
        RECT 121.265 38.385 121.645 38.765 ;
        RECT 121.925 38.385 122.305 38.765 ;
        RECT 122.585 38.385 122.965 38.765 ;
        RECT 121.265 30.305 121.645 30.685 ;
        RECT 121.925 30.305 122.305 30.685 ;
        RECT 122.585 30.305 122.965 30.685 ;
        RECT 121.265 29.645 121.645 30.025 ;
        RECT 121.925 29.645 122.305 30.025 ;
        RECT 122.585 29.645 122.965 30.025 ;
        RECT 121.265 28.985 121.645 29.365 ;
        RECT 121.925 28.985 122.305 29.365 ;
        RECT 122.585 28.985 122.965 29.365 ;
        RECT 132.960 22.205 133.340 22.585 ;
        RECT 133.620 22.205 134.000 22.585 ;
        RECT 134.280 22.205 134.660 22.585 ;
        RECT 132.960 21.545 133.340 21.925 ;
        RECT 133.620 21.545 134.000 21.925 ;
        RECT 134.280 21.545 134.660 21.925 ;
        RECT 132.960 20.885 133.340 21.265 ;
        RECT 133.620 20.885 134.000 21.265 ;
        RECT 134.280 20.885 134.660 21.265 ;
        RECT 94.140 8.770 103.495 9.100 ;
        RECT 94.140 8.750 98.105 8.770 ;
        RECT 72.890 8.090 73.270 8.470 ;
        RECT 87.720 8.090 88.100 8.470 ;
        RECT 72.890 7.430 73.270 7.810 ;
        RECT 87.720 7.430 88.100 7.810 ;
        RECT 72.890 6.770 73.270 7.150 ;
        RECT 87.720 6.770 88.100 7.150 ;
        RECT 70.270 4.690 70.650 5.070 ;
        RECT 76.310 4.720 76.690 5.100 ;
        RECT 76.970 4.720 77.350 5.100 ;
        RECT 77.630 4.720 78.010 5.100 ;
        RECT 82.840 4.690 83.220 5.070 ;
        RECT 83.500 4.690 83.880 5.070 ;
        RECT 84.160 4.690 84.540 5.070 ;
        RECT 91.140 4.720 91.520 5.100 ;
        RECT 91.800 4.720 92.180 5.100 ;
        RECT 92.460 4.720 92.840 5.100 ;
        RECT 97.670 4.690 98.050 5.070 ;
        RECT 98.330 4.690 98.710 5.070 ;
        RECT 98.990 4.690 99.370 5.070 ;
        RECT 101.030 4.690 101.410 5.070 ;
        RECT 101.690 4.690 102.070 5.070 ;
        RECT 102.350 4.690 102.730 5.070 ;
        RECT 53.140 3.420 53.520 3.800 ;
        RECT 69.000 3.770 69.380 4.150 ;
        RECT 52.460 2.580 53.160 2.950 ;
        RECT 53.550 2.760 53.930 3.140 ;
        RECT 55.965 2.950 59.175 3.300 ;
        RECT 52.790 2.305 53.160 2.580 ;
        RECT 55.965 2.305 56.315 2.950 ;
        RECT 60.450 2.760 61.970 3.255 ;
        RECT 63.915 3.125 64.295 3.150 ;
        RECT 62.835 2.795 64.295 3.125 ;
        RECT 60.450 2.600 60.860 2.760 ;
        RECT 52.790 1.955 56.315 2.305 ;
        RECT 56.615 2.250 60.860 2.600 ;
        RECT 46.230 1.555 48.335 1.885 ;
        RECT 61.060 1.885 61.440 1.910 ;
        RECT 62.835 1.885 63.165 2.795 ;
        RECT 63.915 2.770 64.295 2.795 ;
        RECT 71.770 2.950 72.140 4.550 ;
        RECT 72.450 3.420 72.830 3.800 ;
        RECT 71.770 2.580 72.470 2.950 ;
        RECT 72.860 2.760 73.240 3.140 ;
        RECT 75.275 2.950 78.485 3.300 ;
        RECT 72.100 2.305 72.470 2.580 ;
        RECT 75.275 2.305 75.625 2.950 ;
        RECT 79.760 2.760 81.280 3.255 ;
        RECT 83.225 3.125 83.605 3.150 ;
        RECT 82.145 2.795 83.605 3.125 ;
        RECT 79.760 2.600 80.170 2.760 ;
        RECT 72.100 1.955 75.625 2.305 ;
        RECT 75.925 2.250 80.170 2.600 ;
        RECT 61.060 1.555 63.165 1.885 ;
        RECT 80.370 1.885 80.750 1.910 ;
        RECT 82.145 1.885 82.475 2.795 ;
        RECT 83.225 2.770 83.605 2.795 ;
        RECT 86.600 2.950 86.970 4.550 ;
        RECT 103.165 4.150 103.495 8.770 ;
        RECT 114.715 8.750 118.680 9.150 ;
        RECT 136.710 9.150 137.235 59.890 ;
        RECT 138.765 58.745 139.145 59.125 ;
        RECT 138.765 58.085 139.145 58.465 ;
        RECT 138.765 57.425 139.145 57.805 ;
        RECT 138.765 56.765 139.145 57.145 ;
        RECT 138.765 56.105 139.145 56.485 ;
        RECT 138.765 55.445 139.145 55.825 ;
        RECT 138.765 54.785 139.145 55.165 ;
        RECT 138.765 54.125 139.145 54.505 ;
        RECT 138.765 53.465 139.145 53.845 ;
        RECT 138.765 52.805 139.145 53.185 ;
        RECT 138.765 52.145 139.145 52.525 ;
        RECT 138.765 51.485 139.145 51.865 ;
        RECT 138.765 50.825 139.145 51.205 ;
        RECT 138.765 50.165 139.145 50.545 ;
        RECT 140.150 9.150 140.675 59.890 ;
        RECT 149.050 58.745 149.430 59.125 ;
        RECT 149.050 58.085 149.430 58.465 ;
        RECT 149.050 57.425 149.430 57.805 ;
        RECT 149.050 56.765 149.430 57.145 ;
        RECT 149.050 56.105 149.430 56.485 ;
        RECT 149.050 55.445 149.430 55.825 ;
        RECT 149.050 54.785 149.430 55.165 ;
        RECT 149.050 54.125 149.430 54.505 ;
        RECT 149.050 53.465 149.430 53.845 ;
        RECT 149.050 52.805 149.430 53.185 ;
        RECT 149.050 52.145 149.430 52.525 ;
        RECT 149.050 51.485 149.430 51.865 ;
        RECT 149.050 50.825 149.430 51.205 ;
        RECT 149.050 50.165 149.430 50.545 ;
        RECT 143.260 45.105 143.640 45.485 ;
        RECT 143.920 45.105 144.300 45.485 ;
        RECT 144.580 45.105 144.960 45.485 ;
        RECT 143.260 44.445 143.640 44.825 ;
        RECT 143.920 44.445 144.300 44.825 ;
        RECT 144.580 44.445 144.960 44.825 ;
        RECT 143.260 43.785 143.640 44.165 ;
        RECT 143.920 43.785 144.300 44.165 ;
        RECT 144.580 43.785 144.960 44.165 ;
        RECT 153.535 42.405 153.915 42.785 ;
        RECT 154.195 42.405 154.575 42.785 ;
        RECT 154.855 42.405 155.235 42.785 ;
        RECT 153.535 41.745 153.915 42.125 ;
        RECT 154.195 41.745 154.575 42.125 ;
        RECT 154.855 41.745 155.235 42.125 ;
        RECT 153.535 41.085 153.915 41.465 ;
        RECT 154.195 41.085 154.575 41.465 ;
        RECT 154.855 41.085 155.235 41.465 ;
        RECT 153.535 27.605 153.915 27.985 ;
        RECT 154.195 27.605 154.575 27.985 ;
        RECT 154.855 27.605 155.235 27.985 ;
        RECT 153.535 26.945 153.915 27.325 ;
        RECT 154.195 26.945 154.575 27.325 ;
        RECT 154.855 26.945 155.235 27.325 ;
        RECT 153.535 26.285 153.915 26.665 ;
        RECT 154.195 26.285 154.575 26.665 ;
        RECT 154.855 26.285 155.235 26.665 ;
        RECT 143.260 24.905 143.640 25.285 ;
        RECT 143.920 24.905 144.300 25.285 ;
        RECT 144.580 24.905 144.960 25.285 ;
        RECT 143.260 24.245 143.640 24.625 ;
        RECT 143.920 24.245 144.300 24.625 ;
        RECT 144.580 24.245 144.960 24.625 ;
        RECT 143.260 23.585 143.640 23.965 ;
        RECT 143.920 23.585 144.300 23.965 ;
        RECT 144.580 23.585 144.960 23.965 ;
        RECT 136.710 9.100 140.675 9.150 ;
        RECT 157.285 9.150 157.810 59.890 ;
        RECT 159.340 58.745 159.720 59.125 ;
        RECT 159.340 58.085 159.720 58.465 ;
        RECT 159.340 57.425 159.720 57.805 ;
        RECT 159.340 56.765 159.720 57.145 ;
        RECT 159.340 56.105 159.720 56.485 ;
        RECT 159.340 55.445 159.720 55.825 ;
        RECT 159.340 54.785 159.720 55.165 ;
        RECT 159.340 54.125 159.720 54.505 ;
        RECT 159.340 53.465 159.720 53.845 ;
        RECT 159.340 52.805 159.720 53.185 ;
        RECT 159.340 52.145 159.720 52.525 ;
        RECT 159.340 51.485 159.720 51.865 ;
        RECT 159.340 50.825 159.720 51.205 ;
        RECT 159.340 50.165 159.720 50.545 ;
        RECT 160.725 9.150 161.250 59.890 ;
        RECT 169.625 58.745 170.005 59.125 ;
        RECT 171.045 58.745 171.425 59.125 ;
        RECT 169.625 58.085 170.005 58.465 ;
        RECT 171.045 58.085 171.425 58.465 ;
        RECT 169.625 57.425 170.005 57.805 ;
        RECT 171.045 57.425 171.425 57.805 ;
        RECT 169.625 56.765 170.005 57.145 ;
        RECT 171.045 56.765 171.425 57.145 ;
        RECT 169.625 56.105 170.005 56.485 ;
        RECT 171.045 56.105 171.425 56.485 ;
        RECT 169.625 55.445 170.005 55.825 ;
        RECT 171.045 55.445 171.425 55.825 ;
        RECT 169.625 54.785 170.005 55.165 ;
        RECT 171.045 54.785 171.425 55.165 ;
        RECT 169.625 54.125 170.005 54.505 ;
        RECT 171.045 54.125 171.425 54.505 ;
        RECT 169.625 53.465 170.005 53.845 ;
        RECT 171.045 53.465 171.425 53.845 ;
        RECT 169.625 52.805 170.005 53.185 ;
        RECT 171.045 52.805 171.425 53.185 ;
        RECT 169.625 52.145 170.005 52.525 ;
        RECT 171.045 52.145 171.425 52.525 ;
        RECT 169.625 51.485 170.005 51.865 ;
        RECT 171.045 51.485 171.425 51.865 ;
        RECT 169.625 50.825 170.005 51.205 ;
        RECT 171.045 50.825 171.425 51.205 ;
        RECT 169.625 50.165 170.005 50.545 ;
        RECT 171.045 50.165 171.425 50.545 ;
        RECT 175.530 47.805 175.910 48.185 ;
        RECT 176.190 47.805 176.570 48.185 ;
        RECT 176.850 47.805 177.230 48.185 ;
        RECT 175.530 47.145 175.910 47.525 ;
        RECT 176.190 47.145 176.570 47.525 ;
        RECT 176.850 47.145 177.230 47.525 ;
        RECT 175.530 46.485 175.910 46.865 ;
        RECT 176.190 46.485 176.570 46.865 ;
        RECT 176.850 46.485 177.230 46.865 ;
        RECT 163.835 39.705 164.215 40.085 ;
        RECT 164.495 39.705 164.875 40.085 ;
        RECT 165.155 39.705 165.535 40.085 ;
        RECT 163.835 39.045 164.215 39.425 ;
        RECT 164.495 39.045 164.875 39.425 ;
        RECT 165.155 39.045 165.535 39.425 ;
        RECT 163.835 38.385 164.215 38.765 ;
        RECT 164.495 38.385 164.875 38.765 ;
        RECT 165.155 38.385 165.535 38.765 ;
        RECT 163.835 30.305 164.215 30.685 ;
        RECT 164.495 30.305 164.875 30.685 ;
        RECT 165.155 30.305 165.535 30.685 ;
        RECT 163.835 29.645 164.215 30.025 ;
        RECT 164.495 29.645 164.875 30.025 ;
        RECT 165.155 29.645 165.535 30.025 ;
        RECT 163.835 28.985 164.215 29.365 ;
        RECT 164.495 28.985 164.875 29.365 ;
        RECT 165.155 28.985 165.535 29.365 ;
        RECT 175.530 22.205 175.910 22.585 ;
        RECT 176.190 22.205 176.570 22.585 ;
        RECT 176.850 22.205 177.230 22.585 ;
        RECT 175.530 21.545 175.910 21.925 ;
        RECT 176.190 21.545 176.570 21.925 ;
        RECT 176.850 21.545 177.230 21.925 ;
        RECT 175.530 20.885 175.910 21.265 ;
        RECT 176.190 20.885 176.570 21.265 ;
        RECT 176.850 20.885 177.230 21.265 ;
        RECT 136.710 8.770 143.235 9.100 ;
        RECT 136.710 8.750 140.675 8.770 ;
        RECT 107.030 8.090 107.410 8.470 ;
        RECT 121.860 8.090 122.240 8.470 ;
        RECT 107.030 7.430 107.410 7.810 ;
        RECT 121.860 7.430 122.240 7.810 ;
        RECT 107.030 6.770 107.410 7.150 ;
        RECT 121.860 6.770 122.240 7.150 ;
        RECT 104.410 4.690 104.790 5.070 ;
        RECT 110.450 4.720 110.830 5.100 ;
        RECT 111.110 4.720 111.490 5.100 ;
        RECT 111.770 4.720 112.150 5.100 ;
        RECT 116.980 4.690 117.360 5.070 ;
        RECT 117.640 4.690 118.020 5.070 ;
        RECT 118.300 4.690 118.680 5.070 ;
        RECT 125.280 4.720 125.660 5.100 ;
        RECT 125.940 4.720 126.320 5.100 ;
        RECT 126.600 4.720 126.980 5.100 ;
        RECT 131.810 4.690 132.190 5.070 ;
        RECT 132.470 4.690 132.850 5.070 ;
        RECT 133.130 4.690 133.510 5.070 ;
        RECT 135.190 4.690 135.570 5.070 ;
        RECT 136.190 4.690 136.570 5.070 ;
        RECT 136.850 4.690 137.230 5.070 ;
        RECT 137.510 4.690 137.890 5.070 ;
        RECT 138.430 4.690 138.810 5.070 ;
        RECT 139.090 4.690 139.470 5.070 ;
        RECT 139.750 4.690 140.130 5.070 ;
        RECT 140.770 4.690 141.150 5.070 ;
        RECT 141.430 4.690 141.810 5.070 ;
        RECT 142.090 4.690 142.470 5.070 ;
        RECT 87.280 3.420 87.660 3.800 ;
        RECT 103.140 3.770 103.520 4.150 ;
        RECT 86.600 2.580 87.300 2.950 ;
        RECT 87.690 2.760 88.070 3.140 ;
        RECT 90.105 2.950 93.315 3.300 ;
        RECT 86.930 2.305 87.300 2.580 ;
        RECT 90.105 2.305 90.455 2.950 ;
        RECT 94.590 2.760 96.110 3.255 ;
        RECT 98.055 3.125 98.435 3.150 ;
        RECT 96.975 2.795 98.435 3.125 ;
        RECT 94.590 2.600 95.000 2.760 ;
        RECT 86.930 1.955 90.455 2.305 ;
        RECT 90.755 2.250 95.000 2.600 ;
        RECT 80.370 1.555 82.475 1.885 ;
        RECT 95.200 1.885 95.580 1.910 ;
        RECT 96.975 1.885 97.305 2.795 ;
        RECT 98.055 2.770 98.435 2.795 ;
        RECT 105.910 2.950 106.280 4.550 ;
        RECT 106.590 3.420 106.970 3.800 ;
        RECT 105.910 2.580 106.610 2.950 ;
        RECT 107.000 2.760 107.380 3.140 ;
        RECT 109.415 2.950 112.625 3.300 ;
        RECT 106.240 2.305 106.610 2.580 ;
        RECT 109.415 2.305 109.765 2.950 ;
        RECT 113.900 2.760 115.420 3.255 ;
        RECT 117.365 3.125 117.745 3.150 ;
        RECT 116.285 2.795 117.745 3.125 ;
        RECT 113.900 2.600 114.310 2.760 ;
        RECT 106.240 1.955 109.765 2.305 ;
        RECT 110.065 2.250 114.310 2.600 ;
        RECT 95.200 1.555 97.305 1.885 ;
        RECT 114.510 1.885 114.890 1.910 ;
        RECT 116.285 1.885 116.615 2.795 ;
        RECT 117.365 2.770 117.745 2.795 ;
        RECT 120.740 2.950 121.110 4.550 ;
        RECT 142.905 4.150 143.235 8.770 ;
        RECT 157.285 8.750 161.250 9.150 ;
        RECT 179.280 9.150 179.805 59.890 ;
        RECT 181.335 58.745 181.715 59.125 ;
        RECT 181.335 58.085 181.715 58.465 ;
        RECT 181.335 57.425 181.715 57.805 ;
        RECT 181.335 56.765 181.715 57.145 ;
        RECT 181.335 56.105 181.715 56.485 ;
        RECT 181.335 55.445 181.715 55.825 ;
        RECT 181.335 54.785 181.715 55.165 ;
        RECT 181.335 54.125 181.715 54.505 ;
        RECT 181.335 53.465 181.715 53.845 ;
        RECT 181.335 52.805 181.715 53.185 ;
        RECT 181.335 52.145 181.715 52.525 ;
        RECT 181.335 51.485 181.715 51.865 ;
        RECT 181.335 50.825 181.715 51.205 ;
        RECT 181.335 50.165 181.715 50.545 ;
        RECT 182.720 9.150 183.245 59.890 ;
        RECT 191.620 58.745 192.000 59.125 ;
        RECT 191.620 58.085 192.000 58.465 ;
        RECT 191.620 57.425 192.000 57.805 ;
        RECT 191.620 56.765 192.000 57.145 ;
        RECT 191.620 56.105 192.000 56.485 ;
        RECT 191.620 55.445 192.000 55.825 ;
        RECT 191.620 54.785 192.000 55.165 ;
        RECT 191.620 54.125 192.000 54.505 ;
        RECT 191.620 53.465 192.000 53.845 ;
        RECT 191.620 52.805 192.000 53.185 ;
        RECT 191.620 52.145 192.000 52.525 ;
        RECT 191.620 51.485 192.000 51.865 ;
        RECT 191.620 50.825 192.000 51.205 ;
        RECT 191.620 50.165 192.000 50.545 ;
        RECT 185.830 45.105 186.210 45.485 ;
        RECT 186.490 45.105 186.870 45.485 ;
        RECT 187.150 45.105 187.530 45.485 ;
        RECT 185.830 44.445 186.210 44.825 ;
        RECT 186.490 44.445 186.870 44.825 ;
        RECT 187.150 44.445 187.530 44.825 ;
        RECT 185.830 43.785 186.210 44.165 ;
        RECT 186.490 43.785 186.870 44.165 ;
        RECT 187.150 43.785 187.530 44.165 ;
        RECT 196.105 42.405 196.485 42.785 ;
        RECT 196.765 42.405 197.145 42.785 ;
        RECT 197.425 42.405 197.805 42.785 ;
        RECT 196.105 41.745 196.485 42.125 ;
        RECT 196.765 41.745 197.145 42.125 ;
        RECT 197.425 41.745 197.805 42.125 ;
        RECT 196.105 41.085 196.485 41.465 ;
        RECT 196.765 41.085 197.145 41.465 ;
        RECT 197.425 41.085 197.805 41.465 ;
        RECT 196.105 27.605 196.485 27.985 ;
        RECT 196.765 27.605 197.145 27.985 ;
        RECT 197.425 27.605 197.805 27.985 ;
        RECT 196.105 26.945 196.485 27.325 ;
        RECT 196.765 26.945 197.145 27.325 ;
        RECT 197.425 26.945 197.805 27.325 ;
        RECT 196.105 26.285 196.485 26.665 ;
        RECT 196.765 26.285 197.145 26.665 ;
        RECT 197.425 26.285 197.805 26.665 ;
        RECT 185.830 24.905 186.210 25.285 ;
        RECT 186.490 24.905 186.870 25.285 ;
        RECT 187.150 24.905 187.530 25.285 ;
        RECT 185.830 24.245 186.210 24.625 ;
        RECT 186.490 24.245 186.870 24.625 ;
        RECT 187.150 24.245 187.530 24.625 ;
        RECT 185.830 23.585 186.210 23.965 ;
        RECT 186.490 23.585 186.870 23.965 ;
        RECT 187.150 23.585 187.530 23.965 ;
        RECT 179.280 9.100 183.245 9.150 ;
        RECT 199.855 9.150 200.380 59.890 ;
        RECT 201.910 58.745 202.290 59.125 ;
        RECT 201.910 58.085 202.290 58.465 ;
        RECT 201.910 57.425 202.290 57.805 ;
        RECT 201.910 56.765 202.290 57.145 ;
        RECT 201.910 56.105 202.290 56.485 ;
        RECT 201.910 55.445 202.290 55.825 ;
        RECT 201.910 54.785 202.290 55.165 ;
        RECT 201.910 54.125 202.290 54.505 ;
        RECT 201.910 53.465 202.290 53.845 ;
        RECT 201.910 52.805 202.290 53.185 ;
        RECT 201.910 52.145 202.290 52.525 ;
        RECT 201.910 51.485 202.290 51.865 ;
        RECT 201.910 50.825 202.290 51.205 ;
        RECT 201.910 50.165 202.290 50.545 ;
        RECT 203.295 9.150 203.820 59.890 ;
        RECT 212.195 58.745 212.575 59.125 ;
        RECT 213.615 58.745 213.995 59.125 ;
        RECT 212.195 58.085 212.575 58.465 ;
        RECT 213.615 58.085 213.995 58.465 ;
        RECT 212.195 57.425 212.575 57.805 ;
        RECT 213.615 57.425 213.995 57.805 ;
        RECT 212.195 56.765 212.575 57.145 ;
        RECT 213.615 56.765 213.995 57.145 ;
        RECT 212.195 56.105 212.575 56.485 ;
        RECT 213.615 56.105 213.995 56.485 ;
        RECT 212.195 55.445 212.575 55.825 ;
        RECT 213.615 55.445 213.995 55.825 ;
        RECT 212.195 54.785 212.575 55.165 ;
        RECT 213.615 54.785 213.995 55.165 ;
        RECT 212.195 54.125 212.575 54.505 ;
        RECT 213.615 54.125 213.995 54.505 ;
        RECT 212.195 53.465 212.575 53.845 ;
        RECT 213.615 53.465 213.995 53.845 ;
        RECT 212.195 52.805 212.575 53.185 ;
        RECT 213.615 52.805 213.995 53.185 ;
        RECT 212.195 52.145 212.575 52.525 ;
        RECT 213.615 52.145 213.995 52.525 ;
        RECT 212.195 51.485 212.575 51.865 ;
        RECT 213.615 51.485 213.995 51.865 ;
        RECT 212.195 50.825 212.575 51.205 ;
        RECT 213.615 50.825 213.995 51.205 ;
        RECT 212.195 50.165 212.575 50.545 ;
        RECT 213.615 50.165 213.995 50.545 ;
        RECT 218.100 47.805 218.480 48.185 ;
        RECT 218.760 47.805 219.140 48.185 ;
        RECT 219.420 47.805 219.800 48.185 ;
        RECT 218.100 47.145 218.480 47.525 ;
        RECT 218.760 47.145 219.140 47.525 ;
        RECT 219.420 47.145 219.800 47.525 ;
        RECT 218.100 46.485 218.480 46.865 ;
        RECT 218.760 46.485 219.140 46.865 ;
        RECT 219.420 46.485 219.800 46.865 ;
        RECT 206.405 39.705 206.785 40.085 ;
        RECT 207.065 39.705 207.445 40.085 ;
        RECT 207.725 39.705 208.105 40.085 ;
        RECT 206.405 39.045 206.785 39.425 ;
        RECT 207.065 39.045 207.445 39.425 ;
        RECT 207.725 39.045 208.105 39.425 ;
        RECT 206.405 38.385 206.785 38.765 ;
        RECT 207.065 38.385 207.445 38.765 ;
        RECT 207.725 38.385 208.105 38.765 ;
        RECT 206.405 30.305 206.785 30.685 ;
        RECT 207.065 30.305 207.445 30.685 ;
        RECT 207.725 30.305 208.105 30.685 ;
        RECT 206.405 29.645 206.785 30.025 ;
        RECT 207.065 29.645 207.445 30.025 ;
        RECT 207.725 29.645 208.105 30.025 ;
        RECT 206.405 28.985 206.785 29.365 ;
        RECT 207.065 28.985 207.445 29.365 ;
        RECT 207.725 28.985 208.105 29.365 ;
        RECT 218.100 22.205 218.480 22.585 ;
        RECT 218.760 22.205 219.140 22.585 ;
        RECT 219.420 22.205 219.800 22.585 ;
        RECT 218.100 21.545 218.480 21.925 ;
        RECT 218.760 21.545 219.140 21.925 ;
        RECT 219.420 21.545 219.800 21.925 ;
        RECT 218.100 20.885 218.480 21.265 ;
        RECT 218.760 20.885 219.140 21.265 ;
        RECT 219.420 20.885 219.800 21.265 ;
        RECT 179.280 8.770 184.675 9.100 ;
        RECT 179.280 8.750 183.245 8.770 ;
        RECT 144.030 4.690 144.410 5.070 ;
        RECT 144.690 4.690 145.070 5.070 ;
        RECT 145.350 4.690 145.730 5.070 ;
        RECT 146.270 4.690 146.650 5.070 ;
        RECT 146.930 4.690 147.310 5.070 ;
        RECT 147.590 4.690 147.970 5.070 ;
        RECT 148.510 4.690 148.890 5.070 ;
        RECT 149.170 4.690 149.550 5.070 ;
        RECT 149.830 4.690 150.210 5.070 ;
        RECT 150.750 4.690 151.130 5.070 ;
        RECT 151.410 4.690 151.790 5.070 ;
        RECT 152.070 4.690 152.450 5.070 ;
        RECT 152.990 4.690 153.370 5.070 ;
        RECT 153.650 4.690 154.030 5.070 ;
        RECT 154.310 4.690 154.690 5.070 ;
        RECT 155.350 4.690 155.730 5.070 ;
        RECT 156.350 4.690 156.730 5.070 ;
        RECT 157.010 4.690 157.390 5.070 ;
        RECT 157.670 4.690 158.050 5.070 ;
        RECT 158.590 4.690 158.970 5.070 ;
        RECT 159.250 4.690 159.630 5.070 ;
        RECT 159.910 4.690 160.290 5.070 ;
        RECT 160.830 4.690 161.210 5.070 ;
        RECT 161.490 4.690 161.870 5.070 ;
        RECT 162.150 4.690 162.530 5.070 ;
        RECT 163.070 4.690 163.450 5.070 ;
        RECT 163.730 4.690 164.110 5.070 ;
        RECT 164.390 4.690 164.770 5.070 ;
        RECT 165.310 4.690 165.690 5.070 ;
        RECT 165.970 4.690 166.350 5.070 ;
        RECT 166.630 4.690 167.010 5.070 ;
        RECT 167.550 4.690 167.930 5.070 ;
        RECT 168.210 4.690 168.590 5.070 ;
        RECT 168.870 4.690 169.250 5.070 ;
        RECT 169.790 4.690 170.170 5.070 ;
        RECT 170.450 4.690 170.830 5.070 ;
        RECT 171.110 4.690 171.490 5.070 ;
        RECT 172.030 4.690 172.410 5.070 ;
        RECT 172.690 4.690 173.070 5.070 ;
        RECT 173.350 4.690 173.730 5.070 ;
        RECT 174.270 4.690 174.650 5.070 ;
        RECT 174.930 4.690 175.310 5.070 ;
        RECT 175.590 4.690 175.970 5.070 ;
        RECT 176.630 4.690 177.010 5.070 ;
        RECT 177.630 4.690 178.010 5.070 ;
        RECT 178.290 4.690 178.670 5.070 ;
        RECT 178.950 4.690 179.330 5.070 ;
        RECT 179.870 4.690 180.250 5.070 ;
        RECT 180.530 4.690 180.910 5.070 ;
        RECT 181.190 4.690 181.570 5.070 ;
        RECT 182.210 4.690 182.590 5.070 ;
        RECT 182.870 4.690 183.250 5.070 ;
        RECT 183.530 4.690 183.910 5.070 ;
        RECT 184.345 4.150 184.675 8.770 ;
        RECT 199.855 8.750 203.820 9.150 ;
        RECT 221.850 9.150 222.375 59.890 ;
        RECT 223.905 58.745 224.285 59.125 ;
        RECT 223.905 58.085 224.285 58.465 ;
        RECT 223.905 57.425 224.285 57.805 ;
        RECT 223.905 56.765 224.285 57.145 ;
        RECT 223.905 56.105 224.285 56.485 ;
        RECT 223.905 55.445 224.285 55.825 ;
        RECT 223.905 54.785 224.285 55.165 ;
        RECT 223.905 54.125 224.285 54.505 ;
        RECT 223.905 53.465 224.285 53.845 ;
        RECT 223.905 52.805 224.285 53.185 ;
        RECT 223.905 52.145 224.285 52.525 ;
        RECT 223.905 51.485 224.285 51.865 ;
        RECT 223.905 50.825 224.285 51.205 ;
        RECT 223.905 50.165 224.285 50.545 ;
        RECT 225.290 9.150 225.815 59.890 ;
        RECT 234.190 58.745 234.570 59.125 ;
        RECT 234.190 58.085 234.570 58.465 ;
        RECT 234.190 57.425 234.570 57.805 ;
        RECT 234.190 56.765 234.570 57.145 ;
        RECT 234.190 56.105 234.570 56.485 ;
        RECT 234.190 55.445 234.570 55.825 ;
        RECT 234.190 54.785 234.570 55.165 ;
        RECT 234.190 54.125 234.570 54.505 ;
        RECT 234.190 53.465 234.570 53.845 ;
        RECT 234.190 52.805 234.570 53.185 ;
        RECT 234.190 52.145 234.570 52.525 ;
        RECT 234.190 51.485 234.570 51.865 ;
        RECT 234.190 50.825 234.570 51.205 ;
        RECT 234.190 50.165 234.570 50.545 ;
        RECT 228.400 45.105 228.780 45.485 ;
        RECT 229.060 45.105 229.440 45.485 ;
        RECT 229.720 45.105 230.100 45.485 ;
        RECT 228.400 44.445 228.780 44.825 ;
        RECT 229.060 44.445 229.440 44.825 ;
        RECT 229.720 44.445 230.100 44.825 ;
        RECT 228.400 43.785 228.780 44.165 ;
        RECT 229.060 43.785 229.440 44.165 ;
        RECT 229.720 43.785 230.100 44.165 ;
        RECT 238.675 42.405 239.055 42.785 ;
        RECT 239.335 42.405 239.715 42.785 ;
        RECT 239.995 42.405 240.375 42.785 ;
        RECT 238.675 41.745 239.055 42.125 ;
        RECT 239.335 41.745 239.715 42.125 ;
        RECT 239.995 41.745 240.375 42.125 ;
        RECT 238.675 41.085 239.055 41.465 ;
        RECT 239.335 41.085 239.715 41.465 ;
        RECT 239.995 41.085 240.375 41.465 ;
        RECT 238.675 27.605 239.055 27.985 ;
        RECT 239.335 27.605 239.715 27.985 ;
        RECT 239.995 27.605 240.375 27.985 ;
        RECT 238.675 26.945 239.055 27.325 ;
        RECT 239.335 26.945 239.715 27.325 ;
        RECT 239.995 26.945 240.375 27.325 ;
        RECT 238.675 26.285 239.055 26.665 ;
        RECT 239.335 26.285 239.715 26.665 ;
        RECT 239.995 26.285 240.375 26.665 ;
        RECT 228.400 24.905 228.780 25.285 ;
        RECT 229.060 24.905 229.440 25.285 ;
        RECT 229.720 24.905 230.100 25.285 ;
        RECT 228.400 24.245 228.780 24.625 ;
        RECT 229.060 24.245 229.440 24.625 ;
        RECT 229.720 24.245 230.100 24.625 ;
        RECT 228.400 23.585 228.780 23.965 ;
        RECT 229.060 23.585 229.440 23.965 ;
        RECT 229.720 23.585 230.100 23.965 ;
        RECT 221.850 9.100 225.815 9.150 ;
        RECT 242.425 9.150 242.950 59.890 ;
        RECT 244.480 58.745 244.860 59.125 ;
        RECT 244.480 58.085 244.860 58.465 ;
        RECT 244.480 57.425 244.860 57.805 ;
        RECT 244.480 56.765 244.860 57.145 ;
        RECT 244.480 56.105 244.860 56.485 ;
        RECT 244.480 55.445 244.860 55.825 ;
        RECT 244.480 54.785 244.860 55.165 ;
        RECT 244.480 54.125 244.860 54.505 ;
        RECT 244.480 53.465 244.860 53.845 ;
        RECT 244.480 52.805 244.860 53.185 ;
        RECT 244.480 52.145 244.860 52.525 ;
        RECT 244.480 51.485 244.860 51.865 ;
        RECT 244.480 50.825 244.860 51.205 ;
        RECT 244.480 50.165 244.860 50.545 ;
        RECT 245.865 9.150 246.390 59.890 ;
        RECT 254.765 58.745 255.145 59.125 ;
        RECT 256.185 58.745 256.565 59.125 ;
        RECT 254.765 58.085 255.145 58.465 ;
        RECT 256.185 58.085 256.565 58.465 ;
        RECT 254.765 57.425 255.145 57.805 ;
        RECT 256.185 57.425 256.565 57.805 ;
        RECT 254.765 56.765 255.145 57.145 ;
        RECT 256.185 56.765 256.565 57.145 ;
        RECT 254.765 56.105 255.145 56.485 ;
        RECT 256.185 56.105 256.565 56.485 ;
        RECT 254.765 55.445 255.145 55.825 ;
        RECT 256.185 55.445 256.565 55.825 ;
        RECT 254.765 54.785 255.145 55.165 ;
        RECT 256.185 54.785 256.565 55.165 ;
        RECT 254.765 54.125 255.145 54.505 ;
        RECT 256.185 54.125 256.565 54.505 ;
        RECT 254.765 53.465 255.145 53.845 ;
        RECT 256.185 53.465 256.565 53.845 ;
        RECT 254.765 52.805 255.145 53.185 ;
        RECT 256.185 52.805 256.565 53.185 ;
        RECT 254.765 52.145 255.145 52.525 ;
        RECT 256.185 52.145 256.565 52.525 ;
        RECT 254.765 51.485 255.145 51.865 ;
        RECT 256.185 51.485 256.565 51.865 ;
        RECT 254.765 50.825 255.145 51.205 ;
        RECT 256.185 50.825 256.565 51.205 ;
        RECT 254.765 50.165 255.145 50.545 ;
        RECT 256.185 50.165 256.565 50.545 ;
        RECT 260.670 47.805 261.050 48.185 ;
        RECT 261.330 47.805 261.710 48.185 ;
        RECT 261.990 47.805 262.370 48.185 ;
        RECT 260.670 47.145 261.050 47.525 ;
        RECT 261.330 47.145 261.710 47.525 ;
        RECT 261.990 47.145 262.370 47.525 ;
        RECT 260.670 46.485 261.050 46.865 ;
        RECT 261.330 46.485 261.710 46.865 ;
        RECT 261.990 46.485 262.370 46.865 ;
        RECT 248.975 39.705 249.355 40.085 ;
        RECT 249.635 39.705 250.015 40.085 ;
        RECT 250.295 39.705 250.675 40.085 ;
        RECT 248.975 39.045 249.355 39.425 ;
        RECT 249.635 39.045 250.015 39.425 ;
        RECT 250.295 39.045 250.675 39.425 ;
        RECT 248.975 38.385 249.355 38.765 ;
        RECT 249.635 38.385 250.015 38.765 ;
        RECT 250.295 38.385 250.675 38.765 ;
        RECT 248.975 30.305 249.355 30.685 ;
        RECT 249.635 30.305 250.015 30.685 ;
        RECT 250.295 30.305 250.675 30.685 ;
        RECT 248.975 29.645 249.355 30.025 ;
        RECT 249.635 29.645 250.015 30.025 ;
        RECT 250.295 29.645 250.675 30.025 ;
        RECT 248.975 28.985 249.355 29.365 ;
        RECT 249.635 28.985 250.015 29.365 ;
        RECT 250.295 28.985 250.675 29.365 ;
        RECT 260.670 22.205 261.050 22.585 ;
        RECT 261.330 22.205 261.710 22.585 ;
        RECT 261.990 22.205 262.370 22.585 ;
        RECT 260.670 21.545 261.050 21.925 ;
        RECT 261.330 21.545 261.710 21.925 ;
        RECT 261.990 21.545 262.370 21.925 ;
        RECT 260.670 20.885 261.050 21.265 ;
        RECT 261.330 20.885 261.710 21.265 ;
        RECT 261.990 20.885 262.370 21.265 ;
        RECT 221.850 8.770 228.355 9.100 ;
        RECT 221.850 8.750 225.815 8.770 ;
        RECT 185.470 4.690 185.850 5.070 ;
        RECT 186.130 4.690 186.510 5.070 ;
        RECT 186.790 4.690 187.170 5.070 ;
        RECT 187.710 4.690 188.090 5.070 ;
        RECT 188.370 4.690 188.750 5.070 ;
        RECT 189.030 4.690 189.410 5.070 ;
        RECT 189.950 4.690 190.330 5.070 ;
        RECT 190.610 4.690 190.990 5.070 ;
        RECT 191.270 4.690 191.650 5.070 ;
        RECT 192.190 4.690 192.570 5.070 ;
        RECT 192.850 4.690 193.230 5.070 ;
        RECT 193.510 4.690 193.890 5.070 ;
        RECT 194.430 4.690 194.810 5.070 ;
        RECT 195.090 4.690 195.470 5.070 ;
        RECT 195.750 4.690 196.130 5.070 ;
        RECT 196.790 4.690 197.170 5.070 ;
        RECT 197.790 4.690 198.170 5.070 ;
        RECT 198.450 4.690 198.830 5.070 ;
        RECT 199.110 4.690 199.490 5.070 ;
        RECT 200.030 4.690 200.410 5.070 ;
        RECT 200.690 4.690 201.070 5.070 ;
        RECT 201.350 4.690 201.730 5.070 ;
        RECT 202.270 4.690 202.650 5.070 ;
        RECT 202.930 4.690 203.310 5.070 ;
        RECT 203.590 4.690 203.970 5.070 ;
        RECT 204.510 4.690 204.890 5.070 ;
        RECT 205.170 4.690 205.550 5.070 ;
        RECT 205.830 4.690 206.210 5.070 ;
        RECT 206.750 4.690 207.130 5.070 ;
        RECT 207.410 4.690 207.790 5.070 ;
        RECT 208.070 4.690 208.450 5.070 ;
        RECT 208.990 4.690 209.370 5.070 ;
        RECT 209.650 4.690 210.030 5.070 ;
        RECT 210.310 4.690 210.690 5.070 ;
        RECT 211.230 4.690 211.610 5.070 ;
        RECT 211.890 4.690 212.270 5.070 ;
        RECT 212.550 4.690 212.930 5.070 ;
        RECT 213.470 4.690 213.850 5.070 ;
        RECT 214.130 4.690 214.510 5.070 ;
        RECT 214.790 4.690 215.170 5.070 ;
        RECT 215.710 4.690 216.090 5.070 ;
        RECT 216.370 4.690 216.750 5.070 ;
        RECT 217.030 4.690 217.410 5.070 ;
        RECT 218.070 4.690 218.450 5.070 ;
        RECT 219.070 4.690 219.450 5.070 ;
        RECT 219.730 4.690 220.110 5.070 ;
        RECT 220.390 4.690 220.770 5.070 ;
        RECT 221.310 4.690 221.690 5.070 ;
        RECT 221.970 4.690 222.350 5.070 ;
        RECT 222.630 4.690 223.010 5.070 ;
        RECT 223.550 4.690 223.930 5.070 ;
        RECT 224.210 4.690 224.590 5.070 ;
        RECT 224.870 4.690 225.250 5.070 ;
        RECT 225.890 4.690 226.270 5.070 ;
        RECT 226.550 4.690 226.930 5.070 ;
        RECT 227.210 4.690 227.590 5.070 ;
        RECT 228.025 4.150 228.355 8.770 ;
        RECT 242.425 8.750 246.390 9.150 ;
        RECT 264.420 9.150 264.945 59.890 ;
        RECT 266.475 58.745 266.855 59.125 ;
        RECT 266.475 58.085 266.855 58.465 ;
        RECT 266.475 57.425 266.855 57.805 ;
        RECT 266.475 56.765 266.855 57.145 ;
        RECT 266.475 56.105 266.855 56.485 ;
        RECT 266.475 55.445 266.855 55.825 ;
        RECT 266.475 54.785 266.855 55.165 ;
        RECT 266.475 54.125 266.855 54.505 ;
        RECT 266.475 53.465 266.855 53.845 ;
        RECT 266.475 52.805 266.855 53.185 ;
        RECT 266.475 52.145 266.855 52.525 ;
        RECT 266.475 51.485 266.855 51.865 ;
        RECT 266.475 50.825 266.855 51.205 ;
        RECT 266.475 50.165 266.855 50.545 ;
        RECT 267.860 9.150 268.385 59.890 ;
        RECT 276.760 58.745 277.140 59.125 ;
        RECT 276.760 58.085 277.140 58.465 ;
        RECT 276.760 57.425 277.140 57.805 ;
        RECT 276.760 56.765 277.140 57.145 ;
        RECT 276.760 56.105 277.140 56.485 ;
        RECT 276.760 55.445 277.140 55.825 ;
        RECT 276.760 54.785 277.140 55.165 ;
        RECT 276.760 54.125 277.140 54.505 ;
        RECT 276.760 53.465 277.140 53.845 ;
        RECT 276.760 52.805 277.140 53.185 ;
        RECT 276.760 52.145 277.140 52.525 ;
        RECT 276.760 51.485 277.140 51.865 ;
        RECT 276.760 50.825 277.140 51.205 ;
        RECT 276.760 50.165 277.140 50.545 ;
        RECT 270.970 45.105 271.350 45.485 ;
        RECT 271.630 45.105 272.010 45.485 ;
        RECT 272.290 45.105 272.670 45.485 ;
        RECT 270.970 44.445 271.350 44.825 ;
        RECT 271.630 44.445 272.010 44.825 ;
        RECT 272.290 44.445 272.670 44.825 ;
        RECT 270.970 43.785 271.350 44.165 ;
        RECT 271.630 43.785 272.010 44.165 ;
        RECT 272.290 43.785 272.670 44.165 ;
        RECT 281.245 42.405 281.625 42.785 ;
        RECT 281.905 42.405 282.285 42.785 ;
        RECT 282.565 42.405 282.945 42.785 ;
        RECT 281.245 41.745 281.625 42.125 ;
        RECT 281.905 41.745 282.285 42.125 ;
        RECT 282.565 41.745 282.945 42.125 ;
        RECT 281.245 41.085 281.625 41.465 ;
        RECT 281.905 41.085 282.285 41.465 ;
        RECT 282.565 41.085 282.945 41.465 ;
        RECT 281.245 27.605 281.625 27.985 ;
        RECT 281.905 27.605 282.285 27.985 ;
        RECT 282.565 27.605 282.945 27.985 ;
        RECT 281.245 26.945 281.625 27.325 ;
        RECT 281.905 26.945 282.285 27.325 ;
        RECT 282.565 26.945 282.945 27.325 ;
        RECT 281.245 26.285 281.625 26.665 ;
        RECT 281.905 26.285 282.285 26.665 ;
        RECT 282.565 26.285 282.945 26.665 ;
        RECT 270.970 24.905 271.350 25.285 ;
        RECT 271.630 24.905 272.010 25.285 ;
        RECT 272.290 24.905 272.670 25.285 ;
        RECT 270.970 24.245 271.350 24.625 ;
        RECT 271.630 24.245 272.010 24.625 ;
        RECT 272.290 24.245 272.670 24.625 ;
        RECT 270.970 23.585 271.350 23.965 ;
        RECT 271.630 23.585 272.010 23.965 ;
        RECT 272.290 23.585 272.670 23.965 ;
        RECT 264.420 9.100 268.385 9.150 ;
        RECT 284.995 9.150 285.520 59.890 ;
        RECT 287.050 58.745 287.430 59.125 ;
        RECT 287.050 58.085 287.430 58.465 ;
        RECT 287.050 57.425 287.430 57.805 ;
        RECT 287.050 56.765 287.430 57.145 ;
        RECT 287.050 56.105 287.430 56.485 ;
        RECT 287.050 55.445 287.430 55.825 ;
        RECT 287.050 54.785 287.430 55.165 ;
        RECT 287.050 54.125 287.430 54.505 ;
        RECT 287.050 53.465 287.430 53.845 ;
        RECT 287.050 52.805 287.430 53.185 ;
        RECT 287.050 52.145 287.430 52.525 ;
        RECT 287.050 51.485 287.430 51.865 ;
        RECT 287.050 50.825 287.430 51.205 ;
        RECT 287.050 50.165 287.430 50.545 ;
        RECT 288.435 9.150 288.960 59.890 ;
        RECT 297.335 58.745 297.715 59.125 ;
        RECT 298.755 58.745 299.135 59.125 ;
        RECT 297.335 58.085 297.715 58.465 ;
        RECT 298.755 58.085 299.135 58.465 ;
        RECT 297.335 57.425 297.715 57.805 ;
        RECT 298.755 57.425 299.135 57.805 ;
        RECT 297.335 56.765 297.715 57.145 ;
        RECT 298.755 56.765 299.135 57.145 ;
        RECT 297.335 56.105 297.715 56.485 ;
        RECT 298.755 56.105 299.135 56.485 ;
        RECT 297.335 55.445 297.715 55.825 ;
        RECT 298.755 55.445 299.135 55.825 ;
        RECT 297.335 54.785 297.715 55.165 ;
        RECT 298.755 54.785 299.135 55.165 ;
        RECT 297.335 54.125 297.715 54.505 ;
        RECT 298.755 54.125 299.135 54.505 ;
        RECT 297.335 53.465 297.715 53.845 ;
        RECT 298.755 53.465 299.135 53.845 ;
        RECT 297.335 52.805 297.715 53.185 ;
        RECT 298.755 52.805 299.135 53.185 ;
        RECT 297.335 52.145 297.715 52.525 ;
        RECT 298.755 52.145 299.135 52.525 ;
        RECT 297.335 51.485 297.715 51.865 ;
        RECT 298.755 51.485 299.135 51.865 ;
        RECT 297.335 50.825 297.715 51.205 ;
        RECT 298.755 50.825 299.135 51.205 ;
        RECT 297.335 50.165 297.715 50.545 ;
        RECT 298.755 50.165 299.135 50.545 ;
        RECT 303.240 47.805 303.620 48.185 ;
        RECT 303.900 47.805 304.280 48.185 ;
        RECT 304.560 47.805 304.940 48.185 ;
        RECT 303.240 47.145 303.620 47.525 ;
        RECT 303.900 47.145 304.280 47.525 ;
        RECT 304.560 47.145 304.940 47.525 ;
        RECT 303.240 46.485 303.620 46.865 ;
        RECT 303.900 46.485 304.280 46.865 ;
        RECT 304.560 46.485 304.940 46.865 ;
        RECT 291.545 39.705 291.925 40.085 ;
        RECT 292.205 39.705 292.585 40.085 ;
        RECT 292.865 39.705 293.245 40.085 ;
        RECT 291.545 39.045 291.925 39.425 ;
        RECT 292.205 39.045 292.585 39.425 ;
        RECT 292.865 39.045 293.245 39.425 ;
        RECT 291.545 38.385 291.925 38.765 ;
        RECT 292.205 38.385 292.585 38.765 ;
        RECT 292.865 38.385 293.245 38.765 ;
        RECT 291.545 30.305 291.925 30.685 ;
        RECT 292.205 30.305 292.585 30.685 ;
        RECT 292.865 30.305 293.245 30.685 ;
        RECT 291.545 29.645 291.925 30.025 ;
        RECT 292.205 29.645 292.585 30.025 ;
        RECT 292.865 29.645 293.245 30.025 ;
        RECT 291.545 28.985 291.925 29.365 ;
        RECT 292.205 28.985 292.585 29.365 ;
        RECT 292.865 28.985 293.245 29.365 ;
        RECT 303.240 22.205 303.620 22.585 ;
        RECT 303.900 22.205 304.280 22.585 ;
        RECT 304.560 22.205 304.940 22.585 ;
        RECT 303.240 21.545 303.620 21.925 ;
        RECT 303.900 21.545 304.280 21.925 ;
        RECT 304.560 21.545 304.940 21.925 ;
        RECT 303.240 20.885 303.620 21.265 ;
        RECT 303.900 20.885 304.280 21.265 ;
        RECT 304.560 20.885 304.940 21.265 ;
        RECT 264.420 8.770 269.795 9.100 ;
        RECT 264.420 8.750 268.385 8.770 ;
        RECT 229.150 4.690 229.530 5.070 ;
        RECT 229.810 4.690 230.190 5.070 ;
        RECT 230.470 4.690 230.850 5.070 ;
        RECT 231.390 4.690 231.770 5.070 ;
        RECT 232.050 4.690 232.430 5.070 ;
        RECT 232.710 4.690 233.090 5.070 ;
        RECT 233.630 4.690 234.010 5.070 ;
        RECT 234.290 4.690 234.670 5.070 ;
        RECT 234.950 4.690 235.330 5.070 ;
        RECT 235.870 4.690 236.250 5.070 ;
        RECT 236.530 4.690 236.910 5.070 ;
        RECT 237.190 4.690 237.570 5.070 ;
        RECT 238.230 4.690 238.610 5.070 ;
        RECT 239.230 4.690 239.610 5.070 ;
        RECT 239.890 4.690 240.270 5.070 ;
        RECT 240.550 4.690 240.930 5.070 ;
        RECT 241.470 4.690 241.850 5.070 ;
        RECT 242.130 4.690 242.510 5.070 ;
        RECT 242.790 4.690 243.170 5.070 ;
        RECT 243.710 4.690 244.090 5.070 ;
        RECT 244.370 4.690 244.750 5.070 ;
        RECT 245.030 4.690 245.410 5.070 ;
        RECT 245.950 4.690 246.330 5.070 ;
        RECT 246.610 4.690 246.990 5.070 ;
        RECT 247.270 4.690 247.650 5.070 ;
        RECT 248.190 4.690 248.570 5.070 ;
        RECT 248.850 4.690 249.230 5.070 ;
        RECT 249.510 4.690 249.890 5.070 ;
        RECT 250.430 4.690 250.810 5.070 ;
        RECT 251.090 4.690 251.470 5.070 ;
        RECT 251.750 4.690 252.130 5.070 ;
        RECT 252.670 4.690 253.050 5.070 ;
        RECT 253.330 4.690 253.710 5.070 ;
        RECT 253.990 4.690 254.370 5.070 ;
        RECT 254.910 4.690 255.290 5.070 ;
        RECT 255.570 4.690 255.950 5.070 ;
        RECT 256.230 4.690 256.610 5.070 ;
        RECT 257.150 4.690 257.530 5.070 ;
        RECT 257.810 4.690 258.190 5.070 ;
        RECT 258.470 4.690 258.850 5.070 ;
        RECT 259.510 4.690 259.890 5.070 ;
        RECT 260.510 4.690 260.890 5.070 ;
        RECT 261.170 4.690 261.550 5.070 ;
        RECT 261.830 4.690 262.210 5.070 ;
        RECT 262.750 4.690 263.130 5.070 ;
        RECT 263.410 4.690 263.790 5.070 ;
        RECT 264.070 4.690 264.450 5.070 ;
        RECT 264.990 4.690 265.370 5.070 ;
        RECT 265.650 4.690 266.030 5.070 ;
        RECT 266.310 4.690 266.690 5.070 ;
        RECT 267.330 4.690 267.710 5.070 ;
        RECT 267.990 4.690 268.370 5.070 ;
        RECT 268.650 4.690 269.030 5.070 ;
        RECT 269.465 4.150 269.795 8.770 ;
        RECT 284.995 8.750 288.960 9.150 ;
        RECT 306.990 9.150 307.515 59.890 ;
        RECT 309.045 58.745 309.425 59.125 ;
        RECT 309.045 58.085 309.425 58.465 ;
        RECT 309.045 57.425 309.425 57.805 ;
        RECT 309.045 56.765 309.425 57.145 ;
        RECT 309.045 56.105 309.425 56.485 ;
        RECT 309.045 55.445 309.425 55.825 ;
        RECT 309.045 54.785 309.425 55.165 ;
        RECT 309.045 54.125 309.425 54.505 ;
        RECT 309.045 53.465 309.425 53.845 ;
        RECT 309.045 52.805 309.425 53.185 ;
        RECT 309.045 52.145 309.425 52.525 ;
        RECT 309.045 51.485 309.425 51.865 ;
        RECT 309.045 50.825 309.425 51.205 ;
        RECT 309.045 50.165 309.425 50.545 ;
        RECT 310.430 9.150 310.955 59.890 ;
        RECT 319.330 58.745 319.710 59.125 ;
        RECT 319.330 58.085 319.710 58.465 ;
        RECT 319.330 57.425 319.710 57.805 ;
        RECT 319.330 56.765 319.710 57.145 ;
        RECT 319.330 56.105 319.710 56.485 ;
        RECT 319.330 55.445 319.710 55.825 ;
        RECT 319.330 54.785 319.710 55.165 ;
        RECT 319.330 54.125 319.710 54.505 ;
        RECT 319.330 53.465 319.710 53.845 ;
        RECT 319.330 52.805 319.710 53.185 ;
        RECT 319.330 52.145 319.710 52.525 ;
        RECT 319.330 51.485 319.710 51.865 ;
        RECT 319.330 50.825 319.710 51.205 ;
        RECT 319.330 50.165 319.710 50.545 ;
        RECT 313.540 45.105 313.920 45.485 ;
        RECT 314.200 45.105 314.580 45.485 ;
        RECT 314.860 45.105 315.240 45.485 ;
        RECT 313.540 44.445 313.920 44.825 ;
        RECT 314.200 44.445 314.580 44.825 ;
        RECT 314.860 44.445 315.240 44.825 ;
        RECT 313.540 43.785 313.920 44.165 ;
        RECT 314.200 43.785 314.580 44.165 ;
        RECT 314.860 43.785 315.240 44.165 ;
        RECT 323.815 42.405 324.195 42.785 ;
        RECT 324.475 42.405 324.855 42.785 ;
        RECT 325.135 42.405 325.515 42.785 ;
        RECT 323.815 41.745 324.195 42.125 ;
        RECT 324.475 41.745 324.855 42.125 ;
        RECT 325.135 41.745 325.515 42.125 ;
        RECT 323.815 41.085 324.195 41.465 ;
        RECT 324.475 41.085 324.855 41.465 ;
        RECT 325.135 41.085 325.515 41.465 ;
        RECT 323.815 27.605 324.195 27.985 ;
        RECT 324.475 27.605 324.855 27.985 ;
        RECT 325.135 27.605 325.515 27.985 ;
        RECT 323.815 26.945 324.195 27.325 ;
        RECT 324.475 26.945 324.855 27.325 ;
        RECT 325.135 26.945 325.515 27.325 ;
        RECT 323.815 26.285 324.195 26.665 ;
        RECT 324.475 26.285 324.855 26.665 ;
        RECT 325.135 26.285 325.515 26.665 ;
        RECT 313.540 24.905 313.920 25.285 ;
        RECT 314.200 24.905 314.580 25.285 ;
        RECT 314.860 24.905 315.240 25.285 ;
        RECT 313.540 24.245 313.920 24.625 ;
        RECT 314.200 24.245 314.580 24.625 ;
        RECT 314.860 24.245 315.240 24.625 ;
        RECT 313.540 23.585 313.920 23.965 ;
        RECT 314.200 23.585 314.580 23.965 ;
        RECT 314.860 23.585 315.240 23.965 ;
        RECT 306.990 9.100 310.955 9.150 ;
        RECT 327.565 9.150 328.090 59.890 ;
        RECT 329.620 58.745 330.000 59.125 ;
        RECT 329.620 58.085 330.000 58.465 ;
        RECT 329.620 57.425 330.000 57.805 ;
        RECT 329.620 56.765 330.000 57.145 ;
        RECT 329.620 56.105 330.000 56.485 ;
        RECT 329.620 55.445 330.000 55.825 ;
        RECT 329.620 54.785 330.000 55.165 ;
        RECT 329.620 54.125 330.000 54.505 ;
        RECT 329.620 53.465 330.000 53.845 ;
        RECT 329.620 52.805 330.000 53.185 ;
        RECT 329.620 52.145 330.000 52.525 ;
        RECT 329.620 51.485 330.000 51.865 ;
        RECT 329.620 50.825 330.000 51.205 ;
        RECT 329.620 50.165 330.000 50.545 ;
        RECT 331.005 9.150 331.530 59.890 ;
        RECT 339.905 58.745 340.285 59.125 ;
        RECT 341.325 58.745 341.705 59.125 ;
        RECT 339.905 58.085 340.285 58.465 ;
        RECT 341.325 58.085 341.705 58.465 ;
        RECT 339.905 57.425 340.285 57.805 ;
        RECT 341.325 57.425 341.705 57.805 ;
        RECT 339.905 56.765 340.285 57.145 ;
        RECT 341.325 56.765 341.705 57.145 ;
        RECT 339.905 56.105 340.285 56.485 ;
        RECT 341.325 56.105 341.705 56.485 ;
        RECT 339.905 55.445 340.285 55.825 ;
        RECT 341.325 55.445 341.705 55.825 ;
        RECT 339.905 54.785 340.285 55.165 ;
        RECT 341.325 54.785 341.705 55.165 ;
        RECT 339.905 54.125 340.285 54.505 ;
        RECT 341.325 54.125 341.705 54.505 ;
        RECT 339.905 53.465 340.285 53.845 ;
        RECT 341.325 53.465 341.705 53.845 ;
        RECT 339.905 52.805 340.285 53.185 ;
        RECT 341.325 52.805 341.705 53.185 ;
        RECT 339.905 52.145 340.285 52.525 ;
        RECT 341.325 52.145 341.705 52.525 ;
        RECT 339.905 51.485 340.285 51.865 ;
        RECT 341.325 51.485 341.705 51.865 ;
        RECT 339.905 50.825 340.285 51.205 ;
        RECT 341.325 50.825 341.705 51.205 ;
        RECT 339.905 50.165 340.285 50.545 ;
        RECT 341.325 50.165 341.705 50.545 ;
        RECT 345.810 47.805 346.190 48.185 ;
        RECT 346.470 47.805 346.850 48.185 ;
        RECT 347.130 47.805 347.510 48.185 ;
        RECT 345.810 47.145 346.190 47.525 ;
        RECT 346.470 47.145 346.850 47.525 ;
        RECT 347.130 47.145 347.510 47.525 ;
        RECT 345.810 46.485 346.190 46.865 ;
        RECT 346.470 46.485 346.850 46.865 ;
        RECT 347.130 46.485 347.510 46.865 ;
        RECT 334.115 39.705 334.495 40.085 ;
        RECT 334.775 39.705 335.155 40.085 ;
        RECT 335.435 39.705 335.815 40.085 ;
        RECT 334.115 39.045 334.495 39.425 ;
        RECT 334.775 39.045 335.155 39.425 ;
        RECT 335.435 39.045 335.815 39.425 ;
        RECT 334.115 38.385 334.495 38.765 ;
        RECT 334.775 38.385 335.155 38.765 ;
        RECT 335.435 38.385 335.815 38.765 ;
        RECT 334.115 30.305 334.495 30.685 ;
        RECT 334.775 30.305 335.155 30.685 ;
        RECT 335.435 30.305 335.815 30.685 ;
        RECT 334.115 29.645 334.495 30.025 ;
        RECT 334.775 29.645 335.155 30.025 ;
        RECT 335.435 29.645 335.815 30.025 ;
        RECT 334.115 28.985 334.495 29.365 ;
        RECT 334.775 28.985 335.155 29.365 ;
        RECT 335.435 28.985 335.815 29.365 ;
        RECT 345.810 22.205 346.190 22.585 ;
        RECT 346.470 22.205 346.850 22.585 ;
        RECT 347.130 22.205 347.510 22.585 ;
        RECT 345.810 21.545 346.190 21.925 ;
        RECT 346.470 21.545 346.850 21.925 ;
        RECT 347.130 21.545 347.510 21.925 ;
        RECT 345.810 20.885 346.190 21.265 ;
        RECT 346.470 20.885 346.850 21.265 ;
        RECT 347.130 20.885 347.510 21.265 ;
        RECT 306.990 8.770 313.475 9.100 ;
        RECT 306.990 8.750 310.955 8.770 ;
        RECT 270.590 4.690 270.970 5.070 ;
        RECT 271.250 4.690 271.630 5.070 ;
        RECT 271.910 4.690 272.290 5.070 ;
        RECT 272.830 4.690 273.210 5.070 ;
        RECT 273.490 4.690 273.870 5.070 ;
        RECT 274.150 4.690 274.530 5.070 ;
        RECT 275.070 4.690 275.450 5.070 ;
        RECT 275.730 4.690 276.110 5.070 ;
        RECT 276.390 4.690 276.770 5.070 ;
        RECT 277.310 4.690 277.690 5.070 ;
        RECT 277.970 4.690 278.350 5.070 ;
        RECT 278.630 4.690 279.010 5.070 ;
        RECT 279.670 4.690 280.050 5.070 ;
        RECT 280.670 4.690 281.050 5.070 ;
        RECT 281.330 4.690 281.710 5.070 ;
        RECT 281.990 4.690 282.370 5.070 ;
        RECT 282.910 4.690 283.290 5.070 ;
        RECT 283.570 4.690 283.950 5.070 ;
        RECT 284.230 4.690 284.610 5.070 ;
        RECT 285.150 4.690 285.530 5.070 ;
        RECT 285.810 4.690 286.190 5.070 ;
        RECT 286.470 4.690 286.850 5.070 ;
        RECT 287.390 4.690 287.770 5.070 ;
        RECT 288.050 4.690 288.430 5.070 ;
        RECT 288.710 4.690 289.090 5.070 ;
        RECT 289.630 4.690 290.010 5.070 ;
        RECT 290.290 4.690 290.670 5.070 ;
        RECT 290.950 4.690 291.330 5.070 ;
        RECT 291.870 4.690 292.250 5.070 ;
        RECT 292.530 4.690 292.910 5.070 ;
        RECT 293.190 4.690 293.570 5.070 ;
        RECT 294.110 4.690 294.490 5.070 ;
        RECT 294.770 4.690 295.150 5.070 ;
        RECT 295.430 4.690 295.810 5.070 ;
        RECT 296.350 4.690 296.730 5.070 ;
        RECT 297.010 4.690 297.390 5.070 ;
        RECT 297.670 4.690 298.050 5.070 ;
        RECT 298.590 4.690 298.970 5.070 ;
        RECT 299.250 4.690 299.630 5.070 ;
        RECT 299.910 4.690 300.290 5.070 ;
        RECT 300.950 4.690 301.330 5.070 ;
        RECT 301.950 4.690 302.330 5.070 ;
        RECT 302.610 4.690 302.990 5.070 ;
        RECT 303.270 4.690 303.650 5.070 ;
        RECT 304.190 4.690 304.570 5.070 ;
        RECT 304.850 4.690 305.230 5.070 ;
        RECT 305.510 4.690 305.890 5.070 ;
        RECT 306.430 4.690 306.810 5.070 ;
        RECT 307.090 4.690 307.470 5.070 ;
        RECT 307.750 4.690 308.130 5.070 ;
        RECT 308.670 4.690 309.050 5.070 ;
        RECT 309.330 4.690 309.710 5.070 ;
        RECT 309.990 4.690 310.370 5.070 ;
        RECT 311.010 4.690 311.390 5.070 ;
        RECT 311.670 4.690 312.050 5.070 ;
        RECT 312.330 4.690 312.710 5.070 ;
        RECT 313.145 4.150 313.475 8.770 ;
        RECT 327.565 8.750 331.530 9.150 ;
        RECT 349.560 9.150 350.085 59.890 ;
        RECT 351.615 58.745 351.995 59.125 ;
        RECT 351.615 58.085 351.995 58.465 ;
        RECT 351.615 57.425 351.995 57.805 ;
        RECT 351.615 56.765 351.995 57.145 ;
        RECT 351.615 56.105 351.995 56.485 ;
        RECT 351.615 55.445 351.995 55.825 ;
        RECT 351.615 54.785 351.995 55.165 ;
        RECT 351.615 54.125 351.995 54.505 ;
        RECT 351.615 53.465 351.995 53.845 ;
        RECT 351.615 52.805 351.995 53.185 ;
        RECT 351.615 52.145 351.995 52.525 ;
        RECT 351.615 51.485 351.995 51.865 ;
        RECT 351.615 50.825 351.995 51.205 ;
        RECT 351.615 50.165 351.995 50.545 ;
        RECT 353.000 9.150 353.525 59.890 ;
        RECT 361.900 58.745 362.280 59.125 ;
        RECT 361.900 58.085 362.280 58.465 ;
        RECT 361.900 57.425 362.280 57.805 ;
        RECT 361.900 56.765 362.280 57.145 ;
        RECT 361.900 56.105 362.280 56.485 ;
        RECT 361.900 55.445 362.280 55.825 ;
        RECT 361.900 54.785 362.280 55.165 ;
        RECT 361.900 54.125 362.280 54.505 ;
        RECT 361.900 53.465 362.280 53.845 ;
        RECT 361.900 52.805 362.280 53.185 ;
        RECT 361.900 52.145 362.280 52.525 ;
        RECT 361.900 51.485 362.280 51.865 ;
        RECT 361.900 50.825 362.280 51.205 ;
        RECT 361.900 50.165 362.280 50.545 ;
        RECT 356.110 45.105 356.490 45.485 ;
        RECT 356.770 45.105 357.150 45.485 ;
        RECT 357.430 45.105 357.810 45.485 ;
        RECT 356.110 44.445 356.490 44.825 ;
        RECT 356.770 44.445 357.150 44.825 ;
        RECT 357.430 44.445 357.810 44.825 ;
        RECT 356.110 43.785 356.490 44.165 ;
        RECT 356.770 43.785 357.150 44.165 ;
        RECT 357.430 43.785 357.810 44.165 ;
        RECT 366.385 42.405 366.765 42.785 ;
        RECT 367.045 42.405 367.425 42.785 ;
        RECT 367.705 42.405 368.085 42.785 ;
        RECT 366.385 41.745 366.765 42.125 ;
        RECT 367.045 41.745 367.425 42.125 ;
        RECT 367.705 41.745 368.085 42.125 ;
        RECT 366.385 41.085 366.765 41.465 ;
        RECT 367.045 41.085 367.425 41.465 ;
        RECT 367.705 41.085 368.085 41.465 ;
        RECT 366.385 27.605 366.765 27.985 ;
        RECT 367.045 27.605 367.425 27.985 ;
        RECT 367.705 27.605 368.085 27.985 ;
        RECT 366.385 26.945 366.765 27.325 ;
        RECT 367.045 26.945 367.425 27.325 ;
        RECT 367.705 26.945 368.085 27.325 ;
        RECT 366.385 26.285 366.765 26.665 ;
        RECT 367.045 26.285 367.425 26.665 ;
        RECT 367.705 26.285 368.085 26.665 ;
        RECT 356.110 24.905 356.490 25.285 ;
        RECT 356.770 24.905 357.150 25.285 ;
        RECT 357.430 24.905 357.810 25.285 ;
        RECT 356.110 24.245 356.490 24.625 ;
        RECT 356.770 24.245 357.150 24.625 ;
        RECT 357.430 24.245 357.810 24.625 ;
        RECT 356.110 23.585 356.490 23.965 ;
        RECT 356.770 23.585 357.150 23.965 ;
        RECT 357.430 23.585 357.810 23.965 ;
        RECT 349.560 9.100 353.525 9.150 ;
        RECT 370.135 9.150 370.660 59.890 ;
        RECT 372.190 58.745 372.570 59.125 ;
        RECT 372.190 58.085 372.570 58.465 ;
        RECT 372.190 57.425 372.570 57.805 ;
        RECT 372.190 56.765 372.570 57.145 ;
        RECT 372.190 56.105 372.570 56.485 ;
        RECT 372.190 55.445 372.570 55.825 ;
        RECT 372.190 54.785 372.570 55.165 ;
        RECT 372.190 54.125 372.570 54.505 ;
        RECT 372.190 53.465 372.570 53.845 ;
        RECT 372.190 52.805 372.570 53.185 ;
        RECT 372.190 52.145 372.570 52.525 ;
        RECT 372.190 51.485 372.570 51.865 ;
        RECT 372.190 50.825 372.570 51.205 ;
        RECT 372.190 50.165 372.570 50.545 ;
        RECT 373.575 9.150 374.100 59.890 ;
        RECT 382.475 58.745 382.855 59.125 ;
        RECT 383.895 58.745 384.275 59.125 ;
        RECT 382.475 58.085 382.855 58.465 ;
        RECT 383.895 58.085 384.275 58.465 ;
        RECT 382.475 57.425 382.855 57.805 ;
        RECT 383.895 57.425 384.275 57.805 ;
        RECT 382.475 56.765 382.855 57.145 ;
        RECT 383.895 56.765 384.275 57.145 ;
        RECT 382.475 56.105 382.855 56.485 ;
        RECT 383.895 56.105 384.275 56.485 ;
        RECT 382.475 55.445 382.855 55.825 ;
        RECT 383.895 55.445 384.275 55.825 ;
        RECT 382.475 54.785 382.855 55.165 ;
        RECT 383.895 54.785 384.275 55.165 ;
        RECT 382.475 54.125 382.855 54.505 ;
        RECT 383.895 54.125 384.275 54.505 ;
        RECT 382.475 53.465 382.855 53.845 ;
        RECT 383.895 53.465 384.275 53.845 ;
        RECT 382.475 52.805 382.855 53.185 ;
        RECT 383.895 52.805 384.275 53.185 ;
        RECT 382.475 52.145 382.855 52.525 ;
        RECT 383.895 52.145 384.275 52.525 ;
        RECT 382.475 51.485 382.855 51.865 ;
        RECT 383.895 51.485 384.275 51.865 ;
        RECT 382.475 50.825 382.855 51.205 ;
        RECT 383.895 50.825 384.275 51.205 ;
        RECT 382.475 50.165 382.855 50.545 ;
        RECT 383.895 50.165 384.275 50.545 ;
        RECT 388.380 47.805 388.760 48.185 ;
        RECT 389.040 47.805 389.420 48.185 ;
        RECT 389.700 47.805 390.080 48.185 ;
        RECT 388.380 47.145 388.760 47.525 ;
        RECT 389.040 47.145 389.420 47.525 ;
        RECT 389.700 47.145 390.080 47.525 ;
        RECT 388.380 46.485 388.760 46.865 ;
        RECT 389.040 46.485 389.420 46.865 ;
        RECT 389.700 46.485 390.080 46.865 ;
        RECT 376.685 39.705 377.065 40.085 ;
        RECT 377.345 39.705 377.725 40.085 ;
        RECT 378.005 39.705 378.385 40.085 ;
        RECT 376.685 39.045 377.065 39.425 ;
        RECT 377.345 39.045 377.725 39.425 ;
        RECT 378.005 39.045 378.385 39.425 ;
        RECT 376.685 38.385 377.065 38.765 ;
        RECT 377.345 38.385 377.725 38.765 ;
        RECT 378.005 38.385 378.385 38.765 ;
        RECT 376.685 30.305 377.065 30.685 ;
        RECT 377.345 30.305 377.725 30.685 ;
        RECT 378.005 30.305 378.385 30.685 ;
        RECT 376.685 29.645 377.065 30.025 ;
        RECT 377.345 29.645 377.725 30.025 ;
        RECT 378.005 29.645 378.385 30.025 ;
        RECT 376.685 28.985 377.065 29.365 ;
        RECT 377.345 28.985 377.725 29.365 ;
        RECT 378.005 28.985 378.385 29.365 ;
        RECT 388.380 22.205 388.760 22.585 ;
        RECT 389.040 22.205 389.420 22.585 ;
        RECT 389.700 22.205 390.080 22.585 ;
        RECT 388.380 21.545 388.760 21.925 ;
        RECT 389.040 21.545 389.420 21.925 ;
        RECT 389.700 21.545 390.080 21.925 ;
        RECT 388.380 20.885 388.760 21.265 ;
        RECT 389.040 20.885 389.420 21.265 ;
        RECT 389.700 20.885 390.080 21.265 ;
        RECT 349.560 8.770 354.915 9.100 ;
        RECT 349.560 8.750 353.525 8.770 ;
        RECT 314.270 4.690 314.650 5.070 ;
        RECT 314.930 4.690 315.310 5.070 ;
        RECT 315.590 4.690 315.970 5.070 ;
        RECT 316.510 4.690 316.890 5.070 ;
        RECT 317.170 4.690 317.550 5.070 ;
        RECT 317.830 4.690 318.210 5.070 ;
        RECT 318.750 4.690 319.130 5.070 ;
        RECT 319.410 4.690 319.790 5.070 ;
        RECT 320.070 4.690 320.450 5.070 ;
        RECT 321.110 4.690 321.490 5.070 ;
        RECT 322.110 4.690 322.490 5.070 ;
        RECT 322.770 4.690 323.150 5.070 ;
        RECT 323.430 4.690 323.810 5.070 ;
        RECT 324.350 4.690 324.730 5.070 ;
        RECT 325.010 4.690 325.390 5.070 ;
        RECT 325.670 4.690 326.050 5.070 ;
        RECT 326.590 4.690 326.970 5.070 ;
        RECT 327.250 4.690 327.630 5.070 ;
        RECT 327.910 4.690 328.290 5.070 ;
        RECT 328.830 4.690 329.210 5.070 ;
        RECT 329.490 4.690 329.870 5.070 ;
        RECT 330.150 4.690 330.530 5.070 ;
        RECT 331.070 4.690 331.450 5.070 ;
        RECT 331.730 4.690 332.110 5.070 ;
        RECT 332.390 4.690 332.770 5.070 ;
        RECT 333.310 4.690 333.690 5.070 ;
        RECT 333.970 4.690 334.350 5.070 ;
        RECT 334.630 4.690 335.010 5.070 ;
        RECT 335.550 4.690 335.930 5.070 ;
        RECT 336.210 4.690 336.590 5.070 ;
        RECT 336.870 4.690 337.250 5.070 ;
        RECT 337.790 4.690 338.170 5.070 ;
        RECT 338.450 4.690 338.830 5.070 ;
        RECT 339.110 4.690 339.490 5.070 ;
        RECT 340.030 4.690 340.410 5.070 ;
        RECT 340.690 4.690 341.070 5.070 ;
        RECT 341.350 4.690 341.730 5.070 ;
        RECT 342.390 4.690 342.770 5.070 ;
        RECT 343.390 4.690 343.770 5.070 ;
        RECT 344.050 4.690 344.430 5.070 ;
        RECT 344.710 4.690 345.090 5.070 ;
        RECT 345.630 4.690 346.010 5.070 ;
        RECT 346.290 4.690 346.670 5.070 ;
        RECT 346.950 4.690 347.330 5.070 ;
        RECT 347.870 4.690 348.250 5.070 ;
        RECT 348.530 4.690 348.910 5.070 ;
        RECT 349.190 4.690 349.570 5.070 ;
        RECT 350.110 4.690 350.490 5.070 ;
        RECT 350.770 4.690 351.150 5.070 ;
        RECT 351.430 4.690 351.810 5.070 ;
        RECT 352.450 4.690 352.830 5.070 ;
        RECT 353.110 4.690 353.490 5.070 ;
        RECT 353.770 4.690 354.150 5.070 ;
        RECT 354.585 4.150 354.915 8.770 ;
        RECT 370.135 8.750 374.100 9.150 ;
        RECT 392.130 9.150 392.655 59.890 ;
        RECT 394.185 58.745 394.565 59.125 ;
        RECT 394.185 58.085 394.565 58.465 ;
        RECT 394.185 57.425 394.565 57.805 ;
        RECT 394.185 56.765 394.565 57.145 ;
        RECT 394.185 56.105 394.565 56.485 ;
        RECT 394.185 55.445 394.565 55.825 ;
        RECT 394.185 54.785 394.565 55.165 ;
        RECT 394.185 54.125 394.565 54.505 ;
        RECT 394.185 53.465 394.565 53.845 ;
        RECT 394.185 52.805 394.565 53.185 ;
        RECT 394.185 52.145 394.565 52.525 ;
        RECT 394.185 51.485 394.565 51.865 ;
        RECT 394.185 50.825 394.565 51.205 ;
        RECT 394.185 50.165 394.565 50.545 ;
        RECT 395.570 9.150 396.095 59.890 ;
        RECT 404.470 58.745 404.850 59.125 ;
        RECT 404.470 58.085 404.850 58.465 ;
        RECT 404.470 57.425 404.850 57.805 ;
        RECT 404.470 56.765 404.850 57.145 ;
        RECT 404.470 56.105 404.850 56.485 ;
        RECT 404.470 55.445 404.850 55.825 ;
        RECT 404.470 54.785 404.850 55.165 ;
        RECT 404.470 54.125 404.850 54.505 ;
        RECT 404.470 53.465 404.850 53.845 ;
        RECT 404.470 52.805 404.850 53.185 ;
        RECT 404.470 52.145 404.850 52.525 ;
        RECT 404.470 51.485 404.850 51.865 ;
        RECT 404.470 50.825 404.850 51.205 ;
        RECT 404.470 50.165 404.850 50.545 ;
        RECT 398.680 45.105 399.060 45.485 ;
        RECT 399.340 45.105 399.720 45.485 ;
        RECT 400.000 45.105 400.380 45.485 ;
        RECT 398.680 44.445 399.060 44.825 ;
        RECT 399.340 44.445 399.720 44.825 ;
        RECT 400.000 44.445 400.380 44.825 ;
        RECT 398.680 43.785 399.060 44.165 ;
        RECT 399.340 43.785 399.720 44.165 ;
        RECT 400.000 43.785 400.380 44.165 ;
        RECT 408.955 42.405 409.335 42.785 ;
        RECT 409.615 42.405 409.995 42.785 ;
        RECT 410.275 42.405 410.655 42.785 ;
        RECT 408.955 41.745 409.335 42.125 ;
        RECT 409.615 41.745 409.995 42.125 ;
        RECT 410.275 41.745 410.655 42.125 ;
        RECT 408.955 41.085 409.335 41.465 ;
        RECT 409.615 41.085 409.995 41.465 ;
        RECT 410.275 41.085 410.655 41.465 ;
        RECT 408.955 27.605 409.335 27.985 ;
        RECT 409.615 27.605 409.995 27.985 ;
        RECT 410.275 27.605 410.655 27.985 ;
        RECT 408.955 26.945 409.335 27.325 ;
        RECT 409.615 26.945 409.995 27.325 ;
        RECT 410.275 26.945 410.655 27.325 ;
        RECT 408.955 26.285 409.335 26.665 ;
        RECT 409.615 26.285 409.995 26.665 ;
        RECT 410.275 26.285 410.655 26.665 ;
        RECT 398.680 24.905 399.060 25.285 ;
        RECT 399.340 24.905 399.720 25.285 ;
        RECT 400.000 24.905 400.380 25.285 ;
        RECT 398.680 24.245 399.060 24.625 ;
        RECT 399.340 24.245 399.720 24.625 ;
        RECT 400.000 24.245 400.380 24.625 ;
        RECT 398.680 23.585 399.060 23.965 ;
        RECT 399.340 23.585 399.720 23.965 ;
        RECT 400.000 23.585 400.380 23.965 ;
        RECT 392.130 9.100 396.095 9.150 ;
        RECT 412.705 9.150 413.230 59.890 ;
        RECT 414.760 58.745 415.140 59.125 ;
        RECT 414.760 58.085 415.140 58.465 ;
        RECT 414.760 57.425 415.140 57.805 ;
        RECT 414.760 56.765 415.140 57.145 ;
        RECT 414.760 56.105 415.140 56.485 ;
        RECT 414.760 55.445 415.140 55.825 ;
        RECT 414.760 54.785 415.140 55.165 ;
        RECT 414.760 54.125 415.140 54.505 ;
        RECT 414.760 53.465 415.140 53.845 ;
        RECT 414.760 52.805 415.140 53.185 ;
        RECT 414.760 52.145 415.140 52.525 ;
        RECT 414.760 51.485 415.140 51.865 ;
        RECT 414.760 50.825 415.140 51.205 ;
        RECT 414.760 50.165 415.140 50.545 ;
        RECT 416.145 9.150 416.670 59.890 ;
        RECT 425.045 58.745 425.425 59.125 ;
        RECT 426.465 58.745 426.845 59.125 ;
        RECT 425.045 58.085 425.425 58.465 ;
        RECT 426.465 58.085 426.845 58.465 ;
        RECT 425.045 57.425 425.425 57.805 ;
        RECT 426.465 57.425 426.845 57.805 ;
        RECT 425.045 56.765 425.425 57.145 ;
        RECT 426.465 56.765 426.845 57.145 ;
        RECT 425.045 56.105 425.425 56.485 ;
        RECT 426.465 56.105 426.845 56.485 ;
        RECT 425.045 55.445 425.425 55.825 ;
        RECT 426.465 55.445 426.845 55.825 ;
        RECT 425.045 54.785 425.425 55.165 ;
        RECT 426.465 54.785 426.845 55.165 ;
        RECT 425.045 54.125 425.425 54.505 ;
        RECT 426.465 54.125 426.845 54.505 ;
        RECT 425.045 53.465 425.425 53.845 ;
        RECT 426.465 53.465 426.845 53.845 ;
        RECT 425.045 52.805 425.425 53.185 ;
        RECT 426.465 52.805 426.845 53.185 ;
        RECT 425.045 52.145 425.425 52.525 ;
        RECT 426.465 52.145 426.845 52.525 ;
        RECT 425.045 51.485 425.425 51.865 ;
        RECT 426.465 51.485 426.845 51.865 ;
        RECT 425.045 50.825 425.425 51.205 ;
        RECT 426.465 50.825 426.845 51.205 ;
        RECT 425.045 50.165 425.425 50.545 ;
        RECT 426.465 50.165 426.845 50.545 ;
        RECT 430.950 47.805 431.330 48.185 ;
        RECT 431.610 47.805 431.990 48.185 ;
        RECT 432.270 47.805 432.650 48.185 ;
        RECT 430.950 47.145 431.330 47.525 ;
        RECT 431.610 47.145 431.990 47.525 ;
        RECT 432.270 47.145 432.650 47.525 ;
        RECT 430.950 46.485 431.330 46.865 ;
        RECT 431.610 46.485 431.990 46.865 ;
        RECT 432.270 46.485 432.650 46.865 ;
        RECT 419.255 39.705 419.635 40.085 ;
        RECT 419.915 39.705 420.295 40.085 ;
        RECT 420.575 39.705 420.955 40.085 ;
        RECT 419.255 39.045 419.635 39.425 ;
        RECT 419.915 39.045 420.295 39.425 ;
        RECT 420.575 39.045 420.955 39.425 ;
        RECT 419.255 38.385 419.635 38.765 ;
        RECT 419.915 38.385 420.295 38.765 ;
        RECT 420.575 38.385 420.955 38.765 ;
        RECT 419.255 30.305 419.635 30.685 ;
        RECT 419.915 30.305 420.295 30.685 ;
        RECT 420.575 30.305 420.955 30.685 ;
        RECT 419.255 29.645 419.635 30.025 ;
        RECT 419.915 29.645 420.295 30.025 ;
        RECT 420.575 29.645 420.955 30.025 ;
        RECT 419.255 28.985 419.635 29.365 ;
        RECT 419.915 28.985 420.295 29.365 ;
        RECT 420.575 28.985 420.955 29.365 ;
        RECT 430.950 22.205 431.330 22.585 ;
        RECT 431.610 22.205 431.990 22.585 ;
        RECT 432.270 22.205 432.650 22.585 ;
        RECT 430.950 21.545 431.330 21.925 ;
        RECT 431.610 21.545 431.990 21.925 ;
        RECT 432.270 21.545 432.650 21.925 ;
        RECT 430.950 20.885 431.330 21.265 ;
        RECT 431.610 20.885 431.990 21.265 ;
        RECT 432.270 20.885 432.650 21.265 ;
        RECT 392.130 8.770 398.595 9.100 ;
        RECT 392.130 8.750 396.095 8.770 ;
        RECT 355.710 4.690 356.090 5.070 ;
        RECT 356.370 4.690 356.750 5.070 ;
        RECT 357.030 4.690 357.410 5.070 ;
        RECT 357.950 4.690 358.330 5.070 ;
        RECT 358.610 4.690 358.990 5.070 ;
        RECT 359.270 4.690 359.650 5.070 ;
        RECT 360.190 4.690 360.570 5.070 ;
        RECT 360.850 4.690 361.230 5.070 ;
        RECT 361.510 4.690 361.890 5.070 ;
        RECT 362.550 4.690 362.930 5.070 ;
        RECT 363.550 4.690 363.930 5.070 ;
        RECT 364.210 4.690 364.590 5.070 ;
        RECT 364.870 4.690 365.250 5.070 ;
        RECT 365.790 4.690 366.170 5.070 ;
        RECT 366.450 4.690 366.830 5.070 ;
        RECT 367.110 4.690 367.490 5.070 ;
        RECT 368.030 4.690 368.410 5.070 ;
        RECT 368.690 4.690 369.070 5.070 ;
        RECT 369.350 4.690 369.730 5.070 ;
        RECT 370.270 4.690 370.650 5.070 ;
        RECT 370.930 4.690 371.310 5.070 ;
        RECT 371.590 4.690 371.970 5.070 ;
        RECT 372.510 4.690 372.890 5.070 ;
        RECT 373.170 4.690 373.550 5.070 ;
        RECT 373.830 4.690 374.210 5.070 ;
        RECT 374.750 4.690 375.130 5.070 ;
        RECT 375.410 4.690 375.790 5.070 ;
        RECT 376.070 4.690 376.450 5.070 ;
        RECT 376.990 4.690 377.370 5.070 ;
        RECT 377.650 4.690 378.030 5.070 ;
        RECT 378.310 4.690 378.690 5.070 ;
        RECT 379.230 4.690 379.610 5.070 ;
        RECT 379.890 4.690 380.270 5.070 ;
        RECT 380.550 4.690 380.930 5.070 ;
        RECT 381.470 4.690 381.850 5.070 ;
        RECT 382.130 4.690 382.510 5.070 ;
        RECT 382.790 4.690 383.170 5.070 ;
        RECT 383.830 4.690 384.210 5.070 ;
        RECT 384.830 4.690 385.210 5.070 ;
        RECT 385.490 4.690 385.870 5.070 ;
        RECT 386.150 4.690 386.530 5.070 ;
        RECT 387.070 4.690 387.450 5.070 ;
        RECT 387.730 4.690 388.110 5.070 ;
        RECT 388.390 4.690 388.770 5.070 ;
        RECT 389.310 4.690 389.690 5.070 ;
        RECT 389.970 4.690 390.350 5.070 ;
        RECT 390.630 4.690 391.010 5.070 ;
        RECT 391.550 4.690 391.930 5.070 ;
        RECT 392.210 4.690 392.590 5.070 ;
        RECT 392.870 4.690 393.250 5.070 ;
        RECT 393.790 4.690 394.170 5.070 ;
        RECT 394.450 4.690 394.830 5.070 ;
        RECT 395.110 4.690 395.490 5.070 ;
        RECT 396.130 4.690 396.510 5.070 ;
        RECT 396.790 4.690 397.170 5.070 ;
        RECT 397.450 4.690 397.830 5.070 ;
        RECT 398.265 4.150 398.595 8.770 ;
        RECT 412.705 8.750 416.670 9.150 ;
        RECT 434.700 9.150 435.225 59.890 ;
        RECT 436.755 58.745 437.135 59.125 ;
        RECT 436.755 58.085 437.135 58.465 ;
        RECT 436.755 57.425 437.135 57.805 ;
        RECT 436.755 56.765 437.135 57.145 ;
        RECT 436.755 56.105 437.135 56.485 ;
        RECT 436.755 55.445 437.135 55.825 ;
        RECT 436.755 54.785 437.135 55.165 ;
        RECT 436.755 54.125 437.135 54.505 ;
        RECT 436.755 53.465 437.135 53.845 ;
        RECT 436.755 52.805 437.135 53.185 ;
        RECT 436.755 52.145 437.135 52.525 ;
        RECT 436.755 51.485 437.135 51.865 ;
        RECT 436.755 50.825 437.135 51.205 ;
        RECT 436.755 50.165 437.135 50.545 ;
        RECT 438.140 9.150 438.665 59.890 ;
        RECT 447.040 58.745 447.420 59.125 ;
        RECT 447.040 58.085 447.420 58.465 ;
        RECT 447.040 57.425 447.420 57.805 ;
        RECT 447.040 56.765 447.420 57.145 ;
        RECT 447.040 56.105 447.420 56.485 ;
        RECT 447.040 55.445 447.420 55.825 ;
        RECT 447.040 54.785 447.420 55.165 ;
        RECT 447.040 54.125 447.420 54.505 ;
        RECT 447.040 53.465 447.420 53.845 ;
        RECT 447.040 52.805 447.420 53.185 ;
        RECT 447.040 52.145 447.420 52.525 ;
        RECT 447.040 51.485 447.420 51.865 ;
        RECT 447.040 50.825 447.420 51.205 ;
        RECT 447.040 50.165 447.420 50.545 ;
        RECT 441.250 45.105 441.630 45.485 ;
        RECT 441.910 45.105 442.290 45.485 ;
        RECT 442.570 45.105 442.950 45.485 ;
        RECT 441.250 44.445 441.630 44.825 ;
        RECT 441.910 44.445 442.290 44.825 ;
        RECT 442.570 44.445 442.950 44.825 ;
        RECT 441.250 43.785 441.630 44.165 ;
        RECT 441.910 43.785 442.290 44.165 ;
        RECT 442.570 43.785 442.950 44.165 ;
        RECT 451.525 42.405 451.905 42.785 ;
        RECT 452.185 42.405 452.565 42.785 ;
        RECT 452.845 42.405 453.225 42.785 ;
        RECT 451.525 41.745 451.905 42.125 ;
        RECT 452.185 41.745 452.565 42.125 ;
        RECT 452.845 41.745 453.225 42.125 ;
        RECT 451.525 41.085 451.905 41.465 ;
        RECT 452.185 41.085 452.565 41.465 ;
        RECT 452.845 41.085 453.225 41.465 ;
        RECT 451.525 27.605 451.905 27.985 ;
        RECT 452.185 27.605 452.565 27.985 ;
        RECT 452.845 27.605 453.225 27.985 ;
        RECT 451.525 26.945 451.905 27.325 ;
        RECT 452.185 26.945 452.565 27.325 ;
        RECT 452.845 26.945 453.225 27.325 ;
        RECT 451.525 26.285 451.905 26.665 ;
        RECT 452.185 26.285 452.565 26.665 ;
        RECT 452.845 26.285 453.225 26.665 ;
        RECT 441.250 24.905 441.630 25.285 ;
        RECT 441.910 24.905 442.290 25.285 ;
        RECT 442.570 24.905 442.950 25.285 ;
        RECT 441.250 24.245 441.630 24.625 ;
        RECT 441.910 24.245 442.290 24.625 ;
        RECT 442.570 24.245 442.950 24.625 ;
        RECT 441.250 23.585 441.630 23.965 ;
        RECT 441.910 23.585 442.290 23.965 ;
        RECT 442.570 23.585 442.950 23.965 ;
        RECT 434.700 9.100 438.665 9.150 ;
        RECT 455.275 9.150 455.800 59.890 ;
        RECT 457.330 58.745 457.710 59.125 ;
        RECT 457.330 58.085 457.710 58.465 ;
        RECT 457.330 57.425 457.710 57.805 ;
        RECT 457.330 56.765 457.710 57.145 ;
        RECT 457.330 56.105 457.710 56.485 ;
        RECT 457.330 55.445 457.710 55.825 ;
        RECT 457.330 54.785 457.710 55.165 ;
        RECT 457.330 54.125 457.710 54.505 ;
        RECT 457.330 53.465 457.710 53.845 ;
        RECT 457.330 52.805 457.710 53.185 ;
        RECT 457.330 52.145 457.710 52.525 ;
        RECT 457.330 51.485 457.710 51.865 ;
        RECT 457.330 50.825 457.710 51.205 ;
        RECT 457.330 50.165 457.710 50.545 ;
        RECT 458.715 9.150 459.240 59.890 ;
        RECT 467.615 58.745 467.995 59.125 ;
        RECT 469.035 58.745 469.415 59.125 ;
        RECT 467.615 58.085 467.995 58.465 ;
        RECT 469.035 58.085 469.415 58.465 ;
        RECT 467.615 57.425 467.995 57.805 ;
        RECT 469.035 57.425 469.415 57.805 ;
        RECT 467.615 56.765 467.995 57.145 ;
        RECT 469.035 56.765 469.415 57.145 ;
        RECT 467.615 56.105 467.995 56.485 ;
        RECT 469.035 56.105 469.415 56.485 ;
        RECT 467.615 55.445 467.995 55.825 ;
        RECT 469.035 55.445 469.415 55.825 ;
        RECT 467.615 54.785 467.995 55.165 ;
        RECT 469.035 54.785 469.415 55.165 ;
        RECT 467.615 54.125 467.995 54.505 ;
        RECT 469.035 54.125 469.415 54.505 ;
        RECT 467.615 53.465 467.995 53.845 ;
        RECT 469.035 53.465 469.415 53.845 ;
        RECT 467.615 52.805 467.995 53.185 ;
        RECT 469.035 52.805 469.415 53.185 ;
        RECT 467.615 52.145 467.995 52.525 ;
        RECT 469.035 52.145 469.415 52.525 ;
        RECT 467.615 51.485 467.995 51.865 ;
        RECT 469.035 51.485 469.415 51.865 ;
        RECT 467.615 50.825 467.995 51.205 ;
        RECT 469.035 50.825 469.415 51.205 ;
        RECT 467.615 50.165 467.995 50.545 ;
        RECT 469.035 50.165 469.415 50.545 ;
        RECT 473.520 47.805 473.900 48.185 ;
        RECT 474.180 47.805 474.560 48.185 ;
        RECT 474.840 47.805 475.220 48.185 ;
        RECT 473.520 47.145 473.900 47.525 ;
        RECT 474.180 47.145 474.560 47.525 ;
        RECT 474.840 47.145 475.220 47.525 ;
        RECT 473.520 46.485 473.900 46.865 ;
        RECT 474.180 46.485 474.560 46.865 ;
        RECT 474.840 46.485 475.220 46.865 ;
        RECT 461.825 39.705 462.205 40.085 ;
        RECT 462.485 39.705 462.865 40.085 ;
        RECT 463.145 39.705 463.525 40.085 ;
        RECT 461.825 39.045 462.205 39.425 ;
        RECT 462.485 39.045 462.865 39.425 ;
        RECT 463.145 39.045 463.525 39.425 ;
        RECT 461.825 38.385 462.205 38.765 ;
        RECT 462.485 38.385 462.865 38.765 ;
        RECT 463.145 38.385 463.525 38.765 ;
        RECT 461.825 30.305 462.205 30.685 ;
        RECT 462.485 30.305 462.865 30.685 ;
        RECT 463.145 30.305 463.525 30.685 ;
        RECT 461.825 29.645 462.205 30.025 ;
        RECT 462.485 29.645 462.865 30.025 ;
        RECT 463.145 29.645 463.525 30.025 ;
        RECT 461.825 28.985 462.205 29.365 ;
        RECT 462.485 28.985 462.865 29.365 ;
        RECT 463.145 28.985 463.525 29.365 ;
        RECT 473.520 22.205 473.900 22.585 ;
        RECT 474.180 22.205 474.560 22.585 ;
        RECT 474.840 22.205 475.220 22.585 ;
        RECT 473.520 21.545 473.900 21.925 ;
        RECT 474.180 21.545 474.560 21.925 ;
        RECT 474.840 21.545 475.220 21.925 ;
        RECT 473.520 20.885 473.900 21.265 ;
        RECT 474.180 20.885 474.560 21.265 ;
        RECT 474.840 20.885 475.220 21.265 ;
        RECT 434.700 8.770 440.035 9.100 ;
        RECT 434.700 8.750 438.665 8.770 ;
        RECT 399.390 4.690 399.770 5.070 ;
        RECT 400.050 4.690 400.430 5.070 ;
        RECT 400.710 4.690 401.090 5.070 ;
        RECT 401.630 4.690 402.010 5.070 ;
        RECT 402.290 4.690 402.670 5.070 ;
        RECT 402.950 4.690 403.330 5.070 ;
        RECT 403.990 4.690 404.370 5.070 ;
        RECT 404.990 4.690 405.370 5.070 ;
        RECT 405.650 4.690 406.030 5.070 ;
        RECT 406.310 4.690 406.690 5.070 ;
        RECT 407.230 4.690 407.610 5.070 ;
        RECT 407.890 4.690 408.270 5.070 ;
        RECT 408.550 4.690 408.930 5.070 ;
        RECT 409.470 4.690 409.850 5.070 ;
        RECT 410.130 4.690 410.510 5.070 ;
        RECT 410.790 4.690 411.170 5.070 ;
        RECT 411.710 4.690 412.090 5.070 ;
        RECT 412.370 4.690 412.750 5.070 ;
        RECT 413.030 4.690 413.410 5.070 ;
        RECT 413.950 4.690 414.330 5.070 ;
        RECT 414.610 4.690 414.990 5.070 ;
        RECT 415.270 4.690 415.650 5.070 ;
        RECT 416.190 4.690 416.570 5.070 ;
        RECT 416.850 4.690 417.230 5.070 ;
        RECT 417.510 4.690 417.890 5.070 ;
        RECT 418.430 4.690 418.810 5.070 ;
        RECT 419.090 4.690 419.470 5.070 ;
        RECT 419.750 4.690 420.130 5.070 ;
        RECT 420.670 4.690 421.050 5.070 ;
        RECT 421.330 4.690 421.710 5.070 ;
        RECT 421.990 4.690 422.370 5.070 ;
        RECT 422.910 4.690 423.290 5.070 ;
        RECT 423.570 4.690 423.950 5.070 ;
        RECT 424.230 4.690 424.610 5.070 ;
        RECT 425.270 4.690 425.650 5.070 ;
        RECT 426.270 4.690 426.650 5.070 ;
        RECT 426.930 4.690 427.310 5.070 ;
        RECT 427.590 4.690 427.970 5.070 ;
        RECT 428.510 4.690 428.890 5.070 ;
        RECT 429.170 4.690 429.550 5.070 ;
        RECT 429.830 4.690 430.210 5.070 ;
        RECT 430.750 4.690 431.130 5.070 ;
        RECT 431.410 4.690 431.790 5.070 ;
        RECT 432.070 4.690 432.450 5.070 ;
        RECT 432.990 4.690 433.370 5.070 ;
        RECT 433.650 4.690 434.030 5.070 ;
        RECT 434.310 4.690 434.690 5.070 ;
        RECT 435.230 4.690 435.610 5.070 ;
        RECT 435.890 4.690 436.270 5.070 ;
        RECT 436.550 4.690 436.930 5.070 ;
        RECT 437.570 4.690 437.950 5.070 ;
        RECT 438.230 4.690 438.610 5.070 ;
        RECT 438.890 4.690 439.270 5.070 ;
        RECT 439.705 4.150 440.035 8.770 ;
        RECT 455.275 8.750 459.240 9.150 ;
        RECT 477.270 9.150 477.795 59.890 ;
        RECT 479.325 58.745 479.705 59.125 ;
        RECT 479.325 58.085 479.705 58.465 ;
        RECT 479.325 57.425 479.705 57.805 ;
        RECT 479.325 56.765 479.705 57.145 ;
        RECT 479.325 56.105 479.705 56.485 ;
        RECT 479.325 55.445 479.705 55.825 ;
        RECT 479.325 54.785 479.705 55.165 ;
        RECT 479.325 54.125 479.705 54.505 ;
        RECT 479.325 53.465 479.705 53.845 ;
        RECT 479.325 52.805 479.705 53.185 ;
        RECT 479.325 52.145 479.705 52.525 ;
        RECT 479.325 51.485 479.705 51.865 ;
        RECT 479.325 50.825 479.705 51.205 ;
        RECT 479.325 50.165 479.705 50.545 ;
        RECT 480.710 9.150 481.235 59.890 ;
        RECT 489.610 58.745 489.990 59.125 ;
        RECT 489.610 58.085 489.990 58.465 ;
        RECT 489.610 57.425 489.990 57.805 ;
        RECT 489.610 56.765 489.990 57.145 ;
        RECT 489.610 56.105 489.990 56.485 ;
        RECT 489.610 55.445 489.990 55.825 ;
        RECT 489.610 54.785 489.990 55.165 ;
        RECT 489.610 54.125 489.990 54.505 ;
        RECT 489.610 53.465 489.990 53.845 ;
        RECT 489.610 52.805 489.990 53.185 ;
        RECT 489.610 52.145 489.990 52.525 ;
        RECT 489.610 51.485 489.990 51.865 ;
        RECT 489.610 50.825 489.990 51.205 ;
        RECT 489.610 50.165 489.990 50.545 ;
        RECT 483.820 45.105 484.200 45.485 ;
        RECT 484.480 45.105 484.860 45.485 ;
        RECT 485.140 45.105 485.520 45.485 ;
        RECT 483.820 44.445 484.200 44.825 ;
        RECT 484.480 44.445 484.860 44.825 ;
        RECT 485.140 44.445 485.520 44.825 ;
        RECT 483.820 43.785 484.200 44.165 ;
        RECT 484.480 43.785 484.860 44.165 ;
        RECT 485.140 43.785 485.520 44.165 ;
        RECT 494.095 42.405 494.475 42.785 ;
        RECT 494.755 42.405 495.135 42.785 ;
        RECT 495.415 42.405 495.795 42.785 ;
        RECT 494.095 41.745 494.475 42.125 ;
        RECT 494.755 41.745 495.135 42.125 ;
        RECT 495.415 41.745 495.795 42.125 ;
        RECT 494.095 41.085 494.475 41.465 ;
        RECT 494.755 41.085 495.135 41.465 ;
        RECT 495.415 41.085 495.795 41.465 ;
        RECT 494.095 27.605 494.475 27.985 ;
        RECT 494.755 27.605 495.135 27.985 ;
        RECT 495.415 27.605 495.795 27.985 ;
        RECT 494.095 26.945 494.475 27.325 ;
        RECT 494.755 26.945 495.135 27.325 ;
        RECT 495.415 26.945 495.795 27.325 ;
        RECT 494.095 26.285 494.475 26.665 ;
        RECT 494.755 26.285 495.135 26.665 ;
        RECT 495.415 26.285 495.795 26.665 ;
        RECT 483.820 24.905 484.200 25.285 ;
        RECT 484.480 24.905 484.860 25.285 ;
        RECT 485.140 24.905 485.520 25.285 ;
        RECT 483.820 24.245 484.200 24.625 ;
        RECT 484.480 24.245 484.860 24.625 ;
        RECT 485.140 24.245 485.520 24.625 ;
        RECT 483.820 23.585 484.200 23.965 ;
        RECT 484.480 23.585 484.860 23.965 ;
        RECT 485.140 23.585 485.520 23.965 ;
        RECT 477.270 9.100 481.235 9.150 ;
        RECT 497.845 9.150 498.370 59.890 ;
        RECT 499.900 58.745 500.280 59.125 ;
        RECT 499.900 58.085 500.280 58.465 ;
        RECT 499.900 57.425 500.280 57.805 ;
        RECT 499.900 56.765 500.280 57.145 ;
        RECT 499.900 56.105 500.280 56.485 ;
        RECT 499.900 55.445 500.280 55.825 ;
        RECT 499.900 54.785 500.280 55.165 ;
        RECT 499.900 54.125 500.280 54.505 ;
        RECT 499.900 53.465 500.280 53.845 ;
        RECT 499.900 52.805 500.280 53.185 ;
        RECT 499.900 52.145 500.280 52.525 ;
        RECT 499.900 51.485 500.280 51.865 ;
        RECT 499.900 50.825 500.280 51.205 ;
        RECT 499.900 50.165 500.280 50.545 ;
        RECT 501.285 9.150 501.810 59.890 ;
        RECT 510.185 58.745 510.565 59.125 ;
        RECT 511.605 58.745 511.985 59.125 ;
        RECT 510.185 58.085 510.565 58.465 ;
        RECT 511.605 58.085 511.985 58.465 ;
        RECT 510.185 57.425 510.565 57.805 ;
        RECT 511.605 57.425 511.985 57.805 ;
        RECT 510.185 56.765 510.565 57.145 ;
        RECT 511.605 56.765 511.985 57.145 ;
        RECT 510.185 56.105 510.565 56.485 ;
        RECT 511.605 56.105 511.985 56.485 ;
        RECT 510.185 55.445 510.565 55.825 ;
        RECT 511.605 55.445 511.985 55.825 ;
        RECT 510.185 54.785 510.565 55.165 ;
        RECT 511.605 54.785 511.985 55.165 ;
        RECT 510.185 54.125 510.565 54.505 ;
        RECT 511.605 54.125 511.985 54.505 ;
        RECT 510.185 53.465 510.565 53.845 ;
        RECT 511.605 53.465 511.985 53.845 ;
        RECT 510.185 52.805 510.565 53.185 ;
        RECT 511.605 52.805 511.985 53.185 ;
        RECT 510.185 52.145 510.565 52.525 ;
        RECT 511.605 52.145 511.985 52.525 ;
        RECT 510.185 51.485 510.565 51.865 ;
        RECT 511.605 51.485 511.985 51.865 ;
        RECT 510.185 50.825 510.565 51.205 ;
        RECT 511.605 50.825 511.985 51.205 ;
        RECT 510.185 50.165 510.565 50.545 ;
        RECT 511.605 50.165 511.985 50.545 ;
        RECT 516.090 47.805 516.470 48.185 ;
        RECT 516.750 47.805 517.130 48.185 ;
        RECT 517.410 47.805 517.790 48.185 ;
        RECT 516.090 47.145 516.470 47.525 ;
        RECT 516.750 47.145 517.130 47.525 ;
        RECT 517.410 47.145 517.790 47.525 ;
        RECT 516.090 46.485 516.470 46.865 ;
        RECT 516.750 46.485 517.130 46.865 ;
        RECT 517.410 46.485 517.790 46.865 ;
        RECT 504.395 39.705 504.775 40.085 ;
        RECT 505.055 39.705 505.435 40.085 ;
        RECT 505.715 39.705 506.095 40.085 ;
        RECT 504.395 39.045 504.775 39.425 ;
        RECT 505.055 39.045 505.435 39.425 ;
        RECT 505.715 39.045 506.095 39.425 ;
        RECT 504.395 38.385 504.775 38.765 ;
        RECT 505.055 38.385 505.435 38.765 ;
        RECT 505.715 38.385 506.095 38.765 ;
        RECT 504.395 30.305 504.775 30.685 ;
        RECT 505.055 30.305 505.435 30.685 ;
        RECT 505.715 30.305 506.095 30.685 ;
        RECT 504.395 29.645 504.775 30.025 ;
        RECT 505.055 29.645 505.435 30.025 ;
        RECT 505.715 29.645 506.095 30.025 ;
        RECT 504.395 28.985 504.775 29.365 ;
        RECT 505.055 28.985 505.435 29.365 ;
        RECT 505.715 28.985 506.095 29.365 ;
        RECT 516.090 22.205 516.470 22.585 ;
        RECT 516.750 22.205 517.130 22.585 ;
        RECT 517.410 22.205 517.790 22.585 ;
        RECT 516.090 21.545 516.470 21.925 ;
        RECT 516.750 21.545 517.130 21.925 ;
        RECT 517.410 21.545 517.790 21.925 ;
        RECT 516.090 20.885 516.470 21.265 ;
        RECT 516.750 20.885 517.130 21.265 ;
        RECT 517.410 20.885 517.790 21.265 ;
        RECT 477.270 8.770 483.715 9.100 ;
        RECT 477.270 8.750 481.235 8.770 ;
        RECT 440.830 4.690 441.210 5.070 ;
        RECT 441.490 4.690 441.870 5.070 ;
        RECT 442.150 4.690 442.530 5.070 ;
        RECT 443.070 4.690 443.450 5.070 ;
        RECT 443.730 4.690 444.110 5.070 ;
        RECT 444.390 4.690 444.770 5.070 ;
        RECT 445.430 4.690 445.810 5.070 ;
        RECT 446.430 4.690 446.810 5.070 ;
        RECT 447.090 4.690 447.470 5.070 ;
        RECT 447.750 4.690 448.130 5.070 ;
        RECT 448.670 4.690 449.050 5.070 ;
        RECT 449.330 4.690 449.710 5.070 ;
        RECT 449.990 4.690 450.370 5.070 ;
        RECT 450.910 4.690 451.290 5.070 ;
        RECT 451.570 4.690 451.950 5.070 ;
        RECT 452.230 4.690 452.610 5.070 ;
        RECT 453.150 4.690 453.530 5.070 ;
        RECT 453.810 4.690 454.190 5.070 ;
        RECT 454.470 4.690 454.850 5.070 ;
        RECT 455.390 4.690 455.770 5.070 ;
        RECT 456.050 4.690 456.430 5.070 ;
        RECT 456.710 4.690 457.090 5.070 ;
        RECT 457.630 4.690 458.010 5.070 ;
        RECT 458.290 4.690 458.670 5.070 ;
        RECT 458.950 4.690 459.330 5.070 ;
        RECT 459.870 4.690 460.250 5.070 ;
        RECT 460.530 4.690 460.910 5.070 ;
        RECT 461.190 4.690 461.570 5.070 ;
        RECT 462.110 4.690 462.490 5.070 ;
        RECT 462.770 4.690 463.150 5.070 ;
        RECT 463.430 4.690 463.810 5.070 ;
        RECT 464.350 4.690 464.730 5.070 ;
        RECT 465.010 4.690 465.390 5.070 ;
        RECT 465.670 4.690 466.050 5.070 ;
        RECT 466.710 4.690 467.090 5.070 ;
        RECT 467.710 4.690 468.090 5.070 ;
        RECT 468.370 4.690 468.750 5.070 ;
        RECT 469.030 4.690 469.410 5.070 ;
        RECT 469.950 4.690 470.330 5.070 ;
        RECT 470.610 4.690 470.990 5.070 ;
        RECT 471.270 4.690 471.650 5.070 ;
        RECT 472.190 4.690 472.570 5.070 ;
        RECT 472.850 4.690 473.230 5.070 ;
        RECT 473.510 4.690 473.890 5.070 ;
        RECT 474.430 4.690 474.810 5.070 ;
        RECT 475.090 4.690 475.470 5.070 ;
        RECT 475.750 4.690 476.130 5.070 ;
        RECT 476.670 4.690 477.050 5.070 ;
        RECT 477.330 4.690 477.710 5.070 ;
        RECT 477.990 4.690 478.370 5.070 ;
        RECT 478.910 4.690 479.290 5.070 ;
        RECT 479.570 4.690 479.950 5.070 ;
        RECT 480.230 4.690 480.610 5.070 ;
        RECT 481.250 4.690 481.630 5.070 ;
        RECT 481.910 4.690 482.290 5.070 ;
        RECT 482.570 4.690 482.950 5.070 ;
        RECT 483.385 4.150 483.715 8.770 ;
        RECT 497.845 8.750 501.810 9.150 ;
        RECT 519.840 9.150 520.365 59.890 ;
        RECT 521.895 58.745 522.275 59.125 ;
        RECT 521.895 58.085 522.275 58.465 ;
        RECT 521.895 57.425 522.275 57.805 ;
        RECT 521.895 56.765 522.275 57.145 ;
        RECT 521.895 56.105 522.275 56.485 ;
        RECT 521.895 55.445 522.275 55.825 ;
        RECT 521.895 54.785 522.275 55.165 ;
        RECT 521.895 54.125 522.275 54.505 ;
        RECT 521.895 53.465 522.275 53.845 ;
        RECT 521.895 52.805 522.275 53.185 ;
        RECT 521.895 52.145 522.275 52.525 ;
        RECT 521.895 51.485 522.275 51.865 ;
        RECT 521.895 50.825 522.275 51.205 ;
        RECT 521.895 50.165 522.275 50.545 ;
        RECT 523.280 9.150 523.805 59.890 ;
        RECT 532.180 58.745 532.560 59.125 ;
        RECT 532.180 58.085 532.560 58.465 ;
        RECT 532.180 57.425 532.560 57.805 ;
        RECT 532.180 56.765 532.560 57.145 ;
        RECT 532.180 56.105 532.560 56.485 ;
        RECT 532.180 55.445 532.560 55.825 ;
        RECT 532.180 54.785 532.560 55.165 ;
        RECT 532.180 54.125 532.560 54.505 ;
        RECT 532.180 53.465 532.560 53.845 ;
        RECT 532.180 52.805 532.560 53.185 ;
        RECT 532.180 52.145 532.560 52.525 ;
        RECT 532.180 51.485 532.560 51.865 ;
        RECT 532.180 50.825 532.560 51.205 ;
        RECT 532.180 50.165 532.560 50.545 ;
        RECT 526.390 45.105 526.770 45.485 ;
        RECT 527.050 45.105 527.430 45.485 ;
        RECT 527.710 45.105 528.090 45.485 ;
        RECT 526.390 44.445 526.770 44.825 ;
        RECT 527.050 44.445 527.430 44.825 ;
        RECT 527.710 44.445 528.090 44.825 ;
        RECT 526.390 43.785 526.770 44.165 ;
        RECT 527.050 43.785 527.430 44.165 ;
        RECT 527.710 43.785 528.090 44.165 ;
        RECT 536.665 42.405 537.045 42.785 ;
        RECT 537.325 42.405 537.705 42.785 ;
        RECT 537.985 42.405 538.365 42.785 ;
        RECT 536.665 41.745 537.045 42.125 ;
        RECT 537.325 41.745 537.705 42.125 ;
        RECT 537.985 41.745 538.365 42.125 ;
        RECT 536.665 41.085 537.045 41.465 ;
        RECT 537.325 41.085 537.705 41.465 ;
        RECT 537.985 41.085 538.365 41.465 ;
        RECT 536.665 27.605 537.045 27.985 ;
        RECT 537.325 27.605 537.705 27.985 ;
        RECT 537.985 27.605 538.365 27.985 ;
        RECT 536.665 26.945 537.045 27.325 ;
        RECT 537.325 26.945 537.705 27.325 ;
        RECT 537.985 26.945 538.365 27.325 ;
        RECT 536.665 26.285 537.045 26.665 ;
        RECT 537.325 26.285 537.705 26.665 ;
        RECT 537.985 26.285 538.365 26.665 ;
        RECT 526.390 24.905 526.770 25.285 ;
        RECT 527.050 24.905 527.430 25.285 ;
        RECT 527.710 24.905 528.090 25.285 ;
        RECT 526.390 24.245 526.770 24.625 ;
        RECT 527.050 24.245 527.430 24.625 ;
        RECT 527.710 24.245 528.090 24.625 ;
        RECT 526.390 23.585 526.770 23.965 ;
        RECT 527.050 23.585 527.430 23.965 ;
        RECT 527.710 23.585 528.090 23.965 ;
        RECT 519.840 9.100 523.805 9.150 ;
        RECT 540.415 9.150 540.940 59.890 ;
        RECT 542.470 58.745 542.850 59.125 ;
        RECT 542.470 58.085 542.850 58.465 ;
        RECT 542.470 57.425 542.850 57.805 ;
        RECT 542.470 56.765 542.850 57.145 ;
        RECT 542.470 56.105 542.850 56.485 ;
        RECT 542.470 55.445 542.850 55.825 ;
        RECT 542.470 54.785 542.850 55.165 ;
        RECT 542.470 54.125 542.850 54.505 ;
        RECT 542.470 53.465 542.850 53.845 ;
        RECT 542.470 52.805 542.850 53.185 ;
        RECT 542.470 52.145 542.850 52.525 ;
        RECT 542.470 51.485 542.850 51.865 ;
        RECT 542.470 50.825 542.850 51.205 ;
        RECT 542.470 50.165 542.850 50.545 ;
        RECT 543.855 9.150 544.380 59.890 ;
        RECT 552.755 58.745 553.135 59.125 ;
        RECT 554.175 58.745 554.555 59.125 ;
        RECT 552.755 58.085 553.135 58.465 ;
        RECT 554.175 58.085 554.555 58.465 ;
        RECT 552.755 57.425 553.135 57.805 ;
        RECT 554.175 57.425 554.555 57.805 ;
        RECT 552.755 56.765 553.135 57.145 ;
        RECT 554.175 56.765 554.555 57.145 ;
        RECT 552.755 56.105 553.135 56.485 ;
        RECT 554.175 56.105 554.555 56.485 ;
        RECT 552.755 55.445 553.135 55.825 ;
        RECT 554.175 55.445 554.555 55.825 ;
        RECT 552.755 54.785 553.135 55.165 ;
        RECT 554.175 54.785 554.555 55.165 ;
        RECT 552.755 54.125 553.135 54.505 ;
        RECT 554.175 54.125 554.555 54.505 ;
        RECT 552.755 53.465 553.135 53.845 ;
        RECT 554.175 53.465 554.555 53.845 ;
        RECT 552.755 52.805 553.135 53.185 ;
        RECT 554.175 52.805 554.555 53.185 ;
        RECT 552.755 52.145 553.135 52.525 ;
        RECT 554.175 52.145 554.555 52.525 ;
        RECT 552.755 51.485 553.135 51.865 ;
        RECT 554.175 51.485 554.555 51.865 ;
        RECT 552.755 50.825 553.135 51.205 ;
        RECT 554.175 50.825 554.555 51.205 ;
        RECT 552.755 50.165 553.135 50.545 ;
        RECT 554.175 50.165 554.555 50.545 ;
        RECT 558.660 47.805 559.040 48.185 ;
        RECT 559.320 47.805 559.700 48.185 ;
        RECT 559.980 47.805 560.360 48.185 ;
        RECT 558.660 47.145 559.040 47.525 ;
        RECT 559.320 47.145 559.700 47.525 ;
        RECT 559.980 47.145 560.360 47.525 ;
        RECT 558.660 46.485 559.040 46.865 ;
        RECT 559.320 46.485 559.700 46.865 ;
        RECT 559.980 46.485 560.360 46.865 ;
        RECT 546.965 39.705 547.345 40.085 ;
        RECT 547.625 39.705 548.005 40.085 ;
        RECT 548.285 39.705 548.665 40.085 ;
        RECT 546.965 39.045 547.345 39.425 ;
        RECT 547.625 39.045 548.005 39.425 ;
        RECT 548.285 39.045 548.665 39.425 ;
        RECT 546.965 38.385 547.345 38.765 ;
        RECT 547.625 38.385 548.005 38.765 ;
        RECT 548.285 38.385 548.665 38.765 ;
        RECT 546.965 30.305 547.345 30.685 ;
        RECT 547.625 30.305 548.005 30.685 ;
        RECT 548.285 30.305 548.665 30.685 ;
        RECT 546.965 29.645 547.345 30.025 ;
        RECT 547.625 29.645 548.005 30.025 ;
        RECT 548.285 29.645 548.665 30.025 ;
        RECT 546.965 28.985 547.345 29.365 ;
        RECT 547.625 28.985 548.005 29.365 ;
        RECT 548.285 28.985 548.665 29.365 ;
        RECT 558.660 22.205 559.040 22.585 ;
        RECT 559.320 22.205 559.700 22.585 ;
        RECT 559.980 22.205 560.360 22.585 ;
        RECT 558.660 21.545 559.040 21.925 ;
        RECT 559.320 21.545 559.700 21.925 ;
        RECT 559.980 21.545 560.360 21.925 ;
        RECT 558.660 20.885 559.040 21.265 ;
        RECT 559.320 20.885 559.700 21.265 ;
        RECT 559.980 20.885 560.360 21.265 ;
        RECT 519.840 8.770 525.155 9.100 ;
        RECT 519.840 8.750 523.805 8.770 ;
        RECT 484.510 4.690 484.890 5.070 ;
        RECT 485.170 4.690 485.550 5.070 ;
        RECT 485.830 4.690 486.210 5.070 ;
        RECT 486.870 4.690 487.250 5.070 ;
        RECT 487.870 4.690 488.250 5.070 ;
        RECT 488.530 4.690 488.910 5.070 ;
        RECT 489.190 4.690 489.570 5.070 ;
        RECT 490.110 4.690 490.490 5.070 ;
        RECT 490.770 4.690 491.150 5.070 ;
        RECT 491.430 4.690 491.810 5.070 ;
        RECT 492.350 4.690 492.730 5.070 ;
        RECT 493.010 4.690 493.390 5.070 ;
        RECT 493.670 4.690 494.050 5.070 ;
        RECT 494.590 4.690 494.970 5.070 ;
        RECT 495.250 4.690 495.630 5.070 ;
        RECT 495.910 4.690 496.290 5.070 ;
        RECT 496.830 4.690 497.210 5.070 ;
        RECT 497.490 4.690 497.870 5.070 ;
        RECT 498.150 4.690 498.530 5.070 ;
        RECT 499.070 4.690 499.450 5.070 ;
        RECT 499.730 4.690 500.110 5.070 ;
        RECT 500.390 4.690 500.770 5.070 ;
        RECT 501.310 4.690 501.690 5.070 ;
        RECT 501.970 4.690 502.350 5.070 ;
        RECT 502.630 4.690 503.010 5.070 ;
        RECT 503.550 4.690 503.930 5.070 ;
        RECT 504.210 4.690 504.590 5.070 ;
        RECT 504.870 4.690 505.250 5.070 ;
        RECT 505.790 4.690 506.170 5.070 ;
        RECT 506.450 4.690 506.830 5.070 ;
        RECT 507.110 4.690 507.490 5.070 ;
        RECT 508.150 4.690 508.530 5.070 ;
        RECT 509.150 4.690 509.530 5.070 ;
        RECT 509.810 4.690 510.190 5.070 ;
        RECT 510.470 4.690 510.850 5.070 ;
        RECT 511.390 4.690 511.770 5.070 ;
        RECT 512.050 4.690 512.430 5.070 ;
        RECT 512.710 4.690 513.090 5.070 ;
        RECT 513.630 4.690 514.010 5.070 ;
        RECT 514.290 4.690 514.670 5.070 ;
        RECT 514.950 4.690 515.330 5.070 ;
        RECT 515.870 4.690 516.250 5.070 ;
        RECT 516.530 4.690 516.910 5.070 ;
        RECT 517.190 4.690 517.570 5.070 ;
        RECT 518.110 4.690 518.490 5.070 ;
        RECT 518.770 4.690 519.150 5.070 ;
        RECT 519.430 4.690 519.810 5.070 ;
        RECT 520.350 4.690 520.730 5.070 ;
        RECT 521.010 4.690 521.390 5.070 ;
        RECT 521.670 4.690 522.050 5.070 ;
        RECT 522.690 4.690 523.070 5.070 ;
        RECT 523.350 4.690 523.730 5.070 ;
        RECT 524.010 4.690 524.390 5.070 ;
        RECT 524.825 4.150 525.155 8.770 ;
        RECT 540.415 8.750 544.380 9.150 ;
        RECT 562.410 9.150 562.935 59.890 ;
        RECT 564.465 58.745 564.845 59.125 ;
        RECT 564.465 58.085 564.845 58.465 ;
        RECT 564.465 57.425 564.845 57.805 ;
        RECT 564.465 56.765 564.845 57.145 ;
        RECT 564.465 56.105 564.845 56.485 ;
        RECT 564.465 55.445 564.845 55.825 ;
        RECT 564.465 54.785 564.845 55.165 ;
        RECT 564.465 54.125 564.845 54.505 ;
        RECT 564.465 53.465 564.845 53.845 ;
        RECT 564.465 52.805 564.845 53.185 ;
        RECT 564.465 52.145 564.845 52.525 ;
        RECT 564.465 51.485 564.845 51.865 ;
        RECT 564.465 50.825 564.845 51.205 ;
        RECT 564.465 50.165 564.845 50.545 ;
        RECT 565.850 9.150 566.375 59.890 ;
        RECT 574.750 58.745 575.130 59.125 ;
        RECT 574.750 58.085 575.130 58.465 ;
        RECT 574.750 57.425 575.130 57.805 ;
        RECT 574.750 56.765 575.130 57.145 ;
        RECT 574.750 56.105 575.130 56.485 ;
        RECT 574.750 55.445 575.130 55.825 ;
        RECT 574.750 54.785 575.130 55.165 ;
        RECT 574.750 54.125 575.130 54.505 ;
        RECT 574.750 53.465 575.130 53.845 ;
        RECT 574.750 52.805 575.130 53.185 ;
        RECT 574.750 52.145 575.130 52.525 ;
        RECT 574.750 51.485 575.130 51.865 ;
        RECT 574.750 50.825 575.130 51.205 ;
        RECT 574.750 50.165 575.130 50.545 ;
        RECT 568.960 45.105 569.340 45.485 ;
        RECT 569.620 45.105 570.000 45.485 ;
        RECT 570.280 45.105 570.660 45.485 ;
        RECT 568.960 44.445 569.340 44.825 ;
        RECT 569.620 44.445 570.000 44.825 ;
        RECT 570.280 44.445 570.660 44.825 ;
        RECT 568.960 43.785 569.340 44.165 ;
        RECT 569.620 43.785 570.000 44.165 ;
        RECT 570.280 43.785 570.660 44.165 ;
        RECT 579.235 42.405 579.615 42.785 ;
        RECT 579.895 42.405 580.275 42.785 ;
        RECT 580.555 42.405 580.935 42.785 ;
        RECT 579.235 41.745 579.615 42.125 ;
        RECT 579.895 41.745 580.275 42.125 ;
        RECT 580.555 41.745 580.935 42.125 ;
        RECT 579.235 41.085 579.615 41.465 ;
        RECT 579.895 41.085 580.275 41.465 ;
        RECT 580.555 41.085 580.935 41.465 ;
        RECT 579.235 27.605 579.615 27.985 ;
        RECT 579.895 27.605 580.275 27.985 ;
        RECT 580.555 27.605 580.935 27.985 ;
        RECT 579.235 26.945 579.615 27.325 ;
        RECT 579.895 26.945 580.275 27.325 ;
        RECT 580.555 26.945 580.935 27.325 ;
        RECT 579.235 26.285 579.615 26.665 ;
        RECT 579.895 26.285 580.275 26.665 ;
        RECT 580.555 26.285 580.935 26.665 ;
        RECT 568.960 24.905 569.340 25.285 ;
        RECT 569.620 24.905 570.000 25.285 ;
        RECT 570.280 24.905 570.660 25.285 ;
        RECT 568.960 24.245 569.340 24.625 ;
        RECT 569.620 24.245 570.000 24.625 ;
        RECT 570.280 24.245 570.660 24.625 ;
        RECT 568.960 23.585 569.340 23.965 ;
        RECT 569.620 23.585 570.000 23.965 ;
        RECT 570.280 23.585 570.660 23.965 ;
        RECT 562.410 9.100 566.375 9.150 ;
        RECT 582.985 9.150 583.510 59.890 ;
        RECT 585.040 58.745 585.420 59.125 ;
        RECT 585.040 58.085 585.420 58.465 ;
        RECT 585.040 57.425 585.420 57.805 ;
        RECT 585.040 56.765 585.420 57.145 ;
        RECT 585.040 56.105 585.420 56.485 ;
        RECT 585.040 55.445 585.420 55.825 ;
        RECT 585.040 54.785 585.420 55.165 ;
        RECT 585.040 54.125 585.420 54.505 ;
        RECT 585.040 53.465 585.420 53.845 ;
        RECT 585.040 52.805 585.420 53.185 ;
        RECT 585.040 52.145 585.420 52.525 ;
        RECT 585.040 51.485 585.420 51.865 ;
        RECT 585.040 50.825 585.420 51.205 ;
        RECT 585.040 50.165 585.420 50.545 ;
        RECT 586.425 9.150 586.950 59.890 ;
        RECT 595.325 58.745 595.705 59.125 ;
        RECT 596.745 58.745 597.125 59.125 ;
        RECT 595.325 58.085 595.705 58.465 ;
        RECT 596.745 58.085 597.125 58.465 ;
        RECT 595.325 57.425 595.705 57.805 ;
        RECT 596.745 57.425 597.125 57.805 ;
        RECT 595.325 56.765 595.705 57.145 ;
        RECT 596.745 56.765 597.125 57.145 ;
        RECT 595.325 56.105 595.705 56.485 ;
        RECT 596.745 56.105 597.125 56.485 ;
        RECT 595.325 55.445 595.705 55.825 ;
        RECT 596.745 55.445 597.125 55.825 ;
        RECT 595.325 54.785 595.705 55.165 ;
        RECT 596.745 54.785 597.125 55.165 ;
        RECT 595.325 54.125 595.705 54.505 ;
        RECT 596.745 54.125 597.125 54.505 ;
        RECT 595.325 53.465 595.705 53.845 ;
        RECT 596.745 53.465 597.125 53.845 ;
        RECT 595.325 52.805 595.705 53.185 ;
        RECT 596.745 52.805 597.125 53.185 ;
        RECT 595.325 52.145 595.705 52.525 ;
        RECT 596.745 52.145 597.125 52.525 ;
        RECT 595.325 51.485 595.705 51.865 ;
        RECT 596.745 51.485 597.125 51.865 ;
        RECT 595.325 50.825 595.705 51.205 ;
        RECT 596.745 50.825 597.125 51.205 ;
        RECT 595.325 50.165 595.705 50.545 ;
        RECT 596.745 50.165 597.125 50.545 ;
        RECT 601.230 47.805 601.610 48.185 ;
        RECT 601.890 47.805 602.270 48.185 ;
        RECT 602.550 47.805 602.930 48.185 ;
        RECT 601.230 47.145 601.610 47.525 ;
        RECT 601.890 47.145 602.270 47.525 ;
        RECT 602.550 47.145 602.930 47.525 ;
        RECT 601.230 46.485 601.610 46.865 ;
        RECT 601.890 46.485 602.270 46.865 ;
        RECT 602.550 46.485 602.930 46.865 ;
        RECT 589.535 39.705 589.915 40.085 ;
        RECT 590.195 39.705 590.575 40.085 ;
        RECT 590.855 39.705 591.235 40.085 ;
        RECT 589.535 39.045 589.915 39.425 ;
        RECT 590.195 39.045 590.575 39.425 ;
        RECT 590.855 39.045 591.235 39.425 ;
        RECT 589.535 38.385 589.915 38.765 ;
        RECT 590.195 38.385 590.575 38.765 ;
        RECT 590.855 38.385 591.235 38.765 ;
        RECT 589.535 30.305 589.915 30.685 ;
        RECT 590.195 30.305 590.575 30.685 ;
        RECT 590.855 30.305 591.235 30.685 ;
        RECT 589.535 29.645 589.915 30.025 ;
        RECT 590.195 29.645 590.575 30.025 ;
        RECT 590.855 29.645 591.235 30.025 ;
        RECT 589.535 28.985 589.915 29.365 ;
        RECT 590.195 28.985 590.575 29.365 ;
        RECT 590.855 28.985 591.235 29.365 ;
        RECT 601.230 22.205 601.610 22.585 ;
        RECT 601.890 22.205 602.270 22.585 ;
        RECT 602.550 22.205 602.930 22.585 ;
        RECT 601.230 21.545 601.610 21.925 ;
        RECT 601.890 21.545 602.270 21.925 ;
        RECT 602.550 21.545 602.930 21.925 ;
        RECT 601.230 20.885 601.610 21.265 ;
        RECT 601.890 20.885 602.270 21.265 ;
        RECT 602.550 20.885 602.930 21.265 ;
        RECT 562.410 8.770 568.835 9.100 ;
        RECT 562.410 8.750 566.375 8.770 ;
        RECT 525.950 4.690 526.330 5.070 ;
        RECT 526.610 4.690 526.990 5.070 ;
        RECT 527.270 4.690 527.650 5.070 ;
        RECT 528.310 4.690 528.690 5.070 ;
        RECT 529.310 4.690 529.690 5.070 ;
        RECT 529.970 4.690 530.350 5.070 ;
        RECT 530.630 4.690 531.010 5.070 ;
        RECT 531.550 4.690 531.930 5.070 ;
        RECT 532.210 4.690 532.590 5.070 ;
        RECT 532.870 4.690 533.250 5.070 ;
        RECT 533.790 4.690 534.170 5.070 ;
        RECT 534.450 4.690 534.830 5.070 ;
        RECT 535.110 4.690 535.490 5.070 ;
        RECT 536.030 4.690 536.410 5.070 ;
        RECT 536.690 4.690 537.070 5.070 ;
        RECT 537.350 4.690 537.730 5.070 ;
        RECT 538.270 4.690 538.650 5.070 ;
        RECT 538.930 4.690 539.310 5.070 ;
        RECT 539.590 4.690 539.970 5.070 ;
        RECT 540.510 4.690 540.890 5.070 ;
        RECT 541.170 4.690 541.550 5.070 ;
        RECT 541.830 4.690 542.210 5.070 ;
        RECT 542.750 4.690 543.130 5.070 ;
        RECT 543.410 4.690 543.790 5.070 ;
        RECT 544.070 4.690 544.450 5.070 ;
        RECT 544.990 4.690 545.370 5.070 ;
        RECT 545.650 4.690 546.030 5.070 ;
        RECT 546.310 4.690 546.690 5.070 ;
        RECT 547.230 4.690 547.610 5.070 ;
        RECT 547.890 4.690 548.270 5.070 ;
        RECT 548.550 4.690 548.930 5.070 ;
        RECT 549.590 4.690 549.970 5.070 ;
        RECT 550.590 4.690 550.970 5.070 ;
        RECT 551.250 4.690 551.630 5.070 ;
        RECT 551.910 4.690 552.290 5.070 ;
        RECT 552.830 4.690 553.210 5.070 ;
        RECT 553.490 4.690 553.870 5.070 ;
        RECT 554.150 4.690 554.530 5.070 ;
        RECT 555.070 4.690 555.450 5.070 ;
        RECT 555.730 4.690 556.110 5.070 ;
        RECT 556.390 4.690 556.770 5.070 ;
        RECT 557.310 4.690 557.690 5.070 ;
        RECT 557.970 4.690 558.350 5.070 ;
        RECT 558.630 4.690 559.010 5.070 ;
        RECT 559.550 4.690 559.930 5.070 ;
        RECT 560.210 4.690 560.590 5.070 ;
        RECT 560.870 4.690 561.250 5.070 ;
        RECT 561.790 4.690 562.170 5.070 ;
        RECT 562.450 4.690 562.830 5.070 ;
        RECT 563.110 4.690 563.490 5.070 ;
        RECT 564.030 4.690 564.410 5.070 ;
        RECT 564.690 4.690 565.070 5.070 ;
        RECT 565.350 4.690 565.730 5.070 ;
        RECT 566.370 4.690 566.750 5.070 ;
        RECT 567.030 4.690 567.410 5.070 ;
        RECT 567.690 4.690 568.070 5.070 ;
        RECT 568.505 4.150 568.835 8.770 ;
        RECT 582.985 8.750 586.950 9.150 ;
        RECT 604.980 9.150 605.505 59.890 ;
        RECT 607.035 58.745 607.415 59.125 ;
        RECT 607.035 58.085 607.415 58.465 ;
        RECT 607.035 57.425 607.415 57.805 ;
        RECT 607.035 56.765 607.415 57.145 ;
        RECT 607.035 56.105 607.415 56.485 ;
        RECT 607.035 55.445 607.415 55.825 ;
        RECT 607.035 54.785 607.415 55.165 ;
        RECT 607.035 54.125 607.415 54.505 ;
        RECT 607.035 53.465 607.415 53.845 ;
        RECT 607.035 52.805 607.415 53.185 ;
        RECT 607.035 52.145 607.415 52.525 ;
        RECT 607.035 51.485 607.415 51.865 ;
        RECT 607.035 50.825 607.415 51.205 ;
        RECT 607.035 50.165 607.415 50.545 ;
        RECT 608.420 9.150 608.945 59.890 ;
        RECT 617.320 58.745 617.700 59.125 ;
        RECT 617.320 58.085 617.700 58.465 ;
        RECT 617.320 57.425 617.700 57.805 ;
        RECT 617.320 56.765 617.700 57.145 ;
        RECT 617.320 56.105 617.700 56.485 ;
        RECT 617.320 55.445 617.700 55.825 ;
        RECT 617.320 54.785 617.700 55.165 ;
        RECT 617.320 54.125 617.700 54.505 ;
        RECT 617.320 53.465 617.700 53.845 ;
        RECT 617.320 52.805 617.700 53.185 ;
        RECT 617.320 52.145 617.700 52.525 ;
        RECT 617.320 51.485 617.700 51.865 ;
        RECT 617.320 50.825 617.700 51.205 ;
        RECT 617.320 50.165 617.700 50.545 ;
        RECT 611.530 45.105 611.910 45.485 ;
        RECT 612.190 45.105 612.570 45.485 ;
        RECT 612.850 45.105 613.230 45.485 ;
        RECT 611.530 44.445 611.910 44.825 ;
        RECT 612.190 44.445 612.570 44.825 ;
        RECT 612.850 44.445 613.230 44.825 ;
        RECT 611.530 43.785 611.910 44.165 ;
        RECT 612.190 43.785 612.570 44.165 ;
        RECT 612.850 43.785 613.230 44.165 ;
        RECT 621.805 42.405 622.185 42.785 ;
        RECT 622.465 42.405 622.845 42.785 ;
        RECT 623.125 42.405 623.505 42.785 ;
        RECT 621.805 41.745 622.185 42.125 ;
        RECT 622.465 41.745 622.845 42.125 ;
        RECT 623.125 41.745 623.505 42.125 ;
        RECT 621.805 41.085 622.185 41.465 ;
        RECT 622.465 41.085 622.845 41.465 ;
        RECT 623.125 41.085 623.505 41.465 ;
        RECT 621.805 27.605 622.185 27.985 ;
        RECT 622.465 27.605 622.845 27.985 ;
        RECT 623.125 27.605 623.505 27.985 ;
        RECT 621.805 26.945 622.185 27.325 ;
        RECT 622.465 26.945 622.845 27.325 ;
        RECT 623.125 26.945 623.505 27.325 ;
        RECT 621.805 26.285 622.185 26.665 ;
        RECT 622.465 26.285 622.845 26.665 ;
        RECT 623.125 26.285 623.505 26.665 ;
        RECT 611.530 24.905 611.910 25.285 ;
        RECT 612.190 24.905 612.570 25.285 ;
        RECT 612.850 24.905 613.230 25.285 ;
        RECT 611.530 24.245 611.910 24.625 ;
        RECT 612.190 24.245 612.570 24.625 ;
        RECT 612.850 24.245 613.230 24.625 ;
        RECT 611.530 23.585 611.910 23.965 ;
        RECT 612.190 23.585 612.570 23.965 ;
        RECT 612.850 23.585 613.230 23.965 ;
        RECT 604.980 9.100 608.945 9.150 ;
        RECT 625.555 9.150 626.080 59.890 ;
        RECT 627.610 58.745 627.990 59.125 ;
        RECT 627.610 58.085 627.990 58.465 ;
        RECT 627.610 57.425 627.990 57.805 ;
        RECT 627.610 56.765 627.990 57.145 ;
        RECT 627.610 56.105 627.990 56.485 ;
        RECT 627.610 55.445 627.990 55.825 ;
        RECT 627.610 54.785 627.990 55.165 ;
        RECT 627.610 54.125 627.990 54.505 ;
        RECT 627.610 53.465 627.990 53.845 ;
        RECT 627.610 52.805 627.990 53.185 ;
        RECT 627.610 52.145 627.990 52.525 ;
        RECT 627.610 51.485 627.990 51.865 ;
        RECT 627.610 50.825 627.990 51.205 ;
        RECT 627.610 50.165 627.990 50.545 ;
        RECT 628.995 9.150 629.520 59.890 ;
        RECT 637.895 58.745 638.275 59.125 ;
        RECT 639.315 58.745 639.695 59.125 ;
        RECT 637.895 58.085 638.275 58.465 ;
        RECT 639.315 58.085 639.695 58.465 ;
        RECT 637.895 57.425 638.275 57.805 ;
        RECT 639.315 57.425 639.695 57.805 ;
        RECT 637.895 56.765 638.275 57.145 ;
        RECT 639.315 56.765 639.695 57.145 ;
        RECT 637.895 56.105 638.275 56.485 ;
        RECT 639.315 56.105 639.695 56.485 ;
        RECT 637.895 55.445 638.275 55.825 ;
        RECT 639.315 55.445 639.695 55.825 ;
        RECT 637.895 54.785 638.275 55.165 ;
        RECT 639.315 54.785 639.695 55.165 ;
        RECT 637.895 54.125 638.275 54.505 ;
        RECT 639.315 54.125 639.695 54.505 ;
        RECT 637.895 53.465 638.275 53.845 ;
        RECT 639.315 53.465 639.695 53.845 ;
        RECT 637.895 52.805 638.275 53.185 ;
        RECT 639.315 52.805 639.695 53.185 ;
        RECT 637.895 52.145 638.275 52.525 ;
        RECT 639.315 52.145 639.695 52.525 ;
        RECT 637.895 51.485 638.275 51.865 ;
        RECT 639.315 51.485 639.695 51.865 ;
        RECT 637.895 50.825 638.275 51.205 ;
        RECT 639.315 50.825 639.695 51.205 ;
        RECT 637.895 50.165 638.275 50.545 ;
        RECT 639.315 50.165 639.695 50.545 ;
        RECT 643.800 47.805 644.180 48.185 ;
        RECT 644.460 47.805 644.840 48.185 ;
        RECT 645.120 47.805 645.500 48.185 ;
        RECT 643.800 47.145 644.180 47.525 ;
        RECT 644.460 47.145 644.840 47.525 ;
        RECT 645.120 47.145 645.500 47.525 ;
        RECT 643.800 46.485 644.180 46.865 ;
        RECT 644.460 46.485 644.840 46.865 ;
        RECT 645.120 46.485 645.500 46.865 ;
        RECT 632.105 39.705 632.485 40.085 ;
        RECT 632.765 39.705 633.145 40.085 ;
        RECT 633.425 39.705 633.805 40.085 ;
        RECT 632.105 39.045 632.485 39.425 ;
        RECT 632.765 39.045 633.145 39.425 ;
        RECT 633.425 39.045 633.805 39.425 ;
        RECT 632.105 38.385 632.485 38.765 ;
        RECT 632.765 38.385 633.145 38.765 ;
        RECT 633.425 38.385 633.805 38.765 ;
        RECT 632.105 30.305 632.485 30.685 ;
        RECT 632.765 30.305 633.145 30.685 ;
        RECT 633.425 30.305 633.805 30.685 ;
        RECT 632.105 29.645 632.485 30.025 ;
        RECT 632.765 29.645 633.145 30.025 ;
        RECT 633.425 29.645 633.805 30.025 ;
        RECT 632.105 28.985 632.485 29.365 ;
        RECT 632.765 28.985 633.145 29.365 ;
        RECT 633.425 28.985 633.805 29.365 ;
        RECT 643.800 22.205 644.180 22.585 ;
        RECT 644.460 22.205 644.840 22.585 ;
        RECT 645.120 22.205 645.500 22.585 ;
        RECT 643.800 21.545 644.180 21.925 ;
        RECT 644.460 21.545 644.840 21.925 ;
        RECT 645.120 21.545 645.500 21.925 ;
        RECT 643.800 20.885 644.180 21.265 ;
        RECT 644.460 20.885 644.840 21.265 ;
        RECT 645.120 20.885 645.500 21.265 ;
        RECT 604.980 8.770 610.275 9.100 ;
        RECT 604.980 8.750 608.945 8.770 ;
        RECT 569.750 4.690 570.130 5.070 ;
        RECT 570.750 4.690 571.130 5.070 ;
        RECT 571.410 4.690 571.790 5.070 ;
        RECT 572.070 4.690 572.450 5.070 ;
        RECT 572.990 4.690 573.370 5.070 ;
        RECT 573.650 4.690 574.030 5.070 ;
        RECT 574.310 4.690 574.690 5.070 ;
        RECT 575.230 4.690 575.610 5.070 ;
        RECT 575.890 4.690 576.270 5.070 ;
        RECT 576.550 4.690 576.930 5.070 ;
        RECT 577.470 4.690 577.850 5.070 ;
        RECT 578.130 4.690 578.510 5.070 ;
        RECT 578.790 4.690 579.170 5.070 ;
        RECT 579.710 4.690 580.090 5.070 ;
        RECT 580.370 4.690 580.750 5.070 ;
        RECT 581.030 4.690 581.410 5.070 ;
        RECT 581.950 4.690 582.330 5.070 ;
        RECT 582.610 4.690 582.990 5.070 ;
        RECT 583.270 4.690 583.650 5.070 ;
        RECT 584.190 4.690 584.570 5.070 ;
        RECT 584.850 4.690 585.230 5.070 ;
        RECT 585.510 4.690 585.890 5.070 ;
        RECT 586.430 4.690 586.810 5.070 ;
        RECT 587.090 4.690 587.470 5.070 ;
        RECT 587.750 4.690 588.130 5.070 ;
        RECT 588.670 4.690 589.050 5.070 ;
        RECT 589.330 4.690 589.710 5.070 ;
        RECT 589.990 4.690 590.370 5.070 ;
        RECT 591.030 4.690 591.410 5.070 ;
        RECT 592.030 4.690 592.410 5.070 ;
        RECT 592.690 4.690 593.070 5.070 ;
        RECT 593.350 4.690 593.730 5.070 ;
        RECT 594.270 4.690 594.650 5.070 ;
        RECT 594.930 4.690 595.310 5.070 ;
        RECT 595.590 4.690 595.970 5.070 ;
        RECT 596.510 4.690 596.890 5.070 ;
        RECT 597.170 4.690 597.550 5.070 ;
        RECT 597.830 4.690 598.210 5.070 ;
        RECT 598.750 4.690 599.130 5.070 ;
        RECT 599.410 4.690 599.790 5.070 ;
        RECT 600.070 4.690 600.450 5.070 ;
        RECT 600.990 4.690 601.370 5.070 ;
        RECT 601.650 4.690 602.030 5.070 ;
        RECT 602.310 4.690 602.690 5.070 ;
        RECT 603.230 4.690 603.610 5.070 ;
        RECT 603.890 4.690 604.270 5.070 ;
        RECT 604.550 4.690 604.930 5.070 ;
        RECT 605.470 4.690 605.850 5.070 ;
        RECT 606.130 4.690 606.510 5.070 ;
        RECT 606.790 4.690 607.170 5.070 ;
        RECT 607.810 4.690 608.190 5.070 ;
        RECT 608.470 4.690 608.850 5.070 ;
        RECT 609.130 4.690 609.510 5.070 ;
        RECT 609.945 4.150 610.275 8.770 ;
        RECT 625.555 8.750 629.520 9.150 ;
        RECT 647.550 9.150 648.075 59.890 ;
        RECT 649.605 58.745 649.985 59.125 ;
        RECT 649.605 58.085 649.985 58.465 ;
        RECT 649.605 57.425 649.985 57.805 ;
        RECT 649.605 56.765 649.985 57.145 ;
        RECT 649.605 56.105 649.985 56.485 ;
        RECT 649.605 55.445 649.985 55.825 ;
        RECT 649.605 54.785 649.985 55.165 ;
        RECT 649.605 54.125 649.985 54.505 ;
        RECT 649.605 53.465 649.985 53.845 ;
        RECT 649.605 52.805 649.985 53.185 ;
        RECT 649.605 52.145 649.985 52.525 ;
        RECT 649.605 51.485 649.985 51.865 ;
        RECT 649.605 50.825 649.985 51.205 ;
        RECT 649.605 50.165 649.985 50.545 ;
        RECT 650.990 9.150 651.515 59.890 ;
        RECT 659.890 58.745 660.270 59.125 ;
        RECT 659.890 58.085 660.270 58.465 ;
        RECT 659.890 57.425 660.270 57.805 ;
        RECT 659.890 56.765 660.270 57.145 ;
        RECT 659.890 56.105 660.270 56.485 ;
        RECT 659.890 55.445 660.270 55.825 ;
        RECT 659.890 54.785 660.270 55.165 ;
        RECT 659.890 54.125 660.270 54.505 ;
        RECT 659.890 53.465 660.270 53.845 ;
        RECT 659.890 52.805 660.270 53.185 ;
        RECT 659.890 52.145 660.270 52.525 ;
        RECT 659.890 51.485 660.270 51.865 ;
        RECT 659.890 50.825 660.270 51.205 ;
        RECT 659.890 50.165 660.270 50.545 ;
        RECT 654.100 45.105 654.480 45.485 ;
        RECT 654.760 45.105 655.140 45.485 ;
        RECT 655.420 45.105 655.800 45.485 ;
        RECT 654.100 44.445 654.480 44.825 ;
        RECT 654.760 44.445 655.140 44.825 ;
        RECT 655.420 44.445 655.800 44.825 ;
        RECT 654.100 43.785 654.480 44.165 ;
        RECT 654.760 43.785 655.140 44.165 ;
        RECT 655.420 43.785 655.800 44.165 ;
        RECT 664.375 42.405 664.755 42.785 ;
        RECT 665.035 42.405 665.415 42.785 ;
        RECT 665.695 42.405 666.075 42.785 ;
        RECT 664.375 41.745 664.755 42.125 ;
        RECT 665.035 41.745 665.415 42.125 ;
        RECT 665.695 41.745 666.075 42.125 ;
        RECT 664.375 41.085 664.755 41.465 ;
        RECT 665.035 41.085 665.415 41.465 ;
        RECT 665.695 41.085 666.075 41.465 ;
        RECT 664.375 27.605 664.755 27.985 ;
        RECT 665.035 27.605 665.415 27.985 ;
        RECT 665.695 27.605 666.075 27.985 ;
        RECT 664.375 26.945 664.755 27.325 ;
        RECT 665.035 26.945 665.415 27.325 ;
        RECT 665.695 26.945 666.075 27.325 ;
        RECT 664.375 26.285 664.755 26.665 ;
        RECT 665.035 26.285 665.415 26.665 ;
        RECT 665.695 26.285 666.075 26.665 ;
        RECT 654.100 24.905 654.480 25.285 ;
        RECT 654.760 24.905 655.140 25.285 ;
        RECT 655.420 24.905 655.800 25.285 ;
        RECT 654.100 24.245 654.480 24.625 ;
        RECT 654.760 24.245 655.140 24.625 ;
        RECT 655.420 24.245 655.800 24.625 ;
        RECT 654.100 23.585 654.480 23.965 ;
        RECT 654.760 23.585 655.140 23.965 ;
        RECT 655.420 23.585 655.800 23.965 ;
        RECT 647.550 9.100 651.515 9.150 ;
        RECT 668.125 9.150 668.650 59.890 ;
        RECT 670.180 58.745 670.560 59.125 ;
        RECT 670.180 58.085 670.560 58.465 ;
        RECT 670.180 57.425 670.560 57.805 ;
        RECT 670.180 56.765 670.560 57.145 ;
        RECT 670.180 56.105 670.560 56.485 ;
        RECT 670.180 55.445 670.560 55.825 ;
        RECT 670.180 54.785 670.560 55.165 ;
        RECT 670.180 54.125 670.560 54.505 ;
        RECT 670.180 53.465 670.560 53.845 ;
        RECT 670.180 52.805 670.560 53.185 ;
        RECT 670.180 52.145 670.560 52.525 ;
        RECT 670.180 51.485 670.560 51.865 ;
        RECT 670.180 50.825 670.560 51.205 ;
        RECT 670.180 50.165 670.560 50.545 ;
        RECT 671.565 9.150 672.090 59.890 ;
        RECT 680.465 58.745 680.845 59.125 ;
        RECT 680.465 58.085 680.845 58.465 ;
        RECT 680.465 57.425 680.845 57.805 ;
        RECT 680.465 56.765 680.845 57.145 ;
        RECT 680.465 56.105 680.845 56.485 ;
        RECT 680.465 55.445 680.845 55.825 ;
        RECT 680.465 54.785 680.845 55.165 ;
        RECT 682.310 55.115 682.690 55.495 ;
        RECT 684.095 55.115 684.475 55.495 ;
        RECT 686.950 55.115 687.330 55.495 ;
        RECT 688.735 55.115 689.115 55.495 ;
        RECT 691.590 55.115 691.970 55.495 ;
        RECT 693.375 55.115 693.755 55.495 ;
        RECT 696.230 55.115 696.610 55.495 ;
        RECT 698.015 55.115 698.395 55.495 ;
        RECT 700.870 55.115 701.250 55.495 ;
        RECT 702.655 55.115 703.035 55.495 ;
        RECT 705.510 55.115 705.890 55.495 ;
        RECT 707.295 55.115 707.675 55.495 ;
        RECT 710.150 55.115 710.530 55.495 ;
        RECT 711.935 55.115 712.315 55.495 ;
        RECT 714.790 55.115 715.170 55.495 ;
        RECT 716.575 55.115 716.955 55.495 ;
        RECT 680.465 54.125 680.845 54.505 ;
        RECT 682.310 54.455 682.690 54.835 ;
        RECT 684.095 54.455 684.475 54.835 ;
        RECT 686.950 54.455 687.330 54.835 ;
        RECT 688.735 54.455 689.115 54.835 ;
        RECT 691.590 54.455 691.970 54.835 ;
        RECT 693.375 54.455 693.755 54.835 ;
        RECT 696.230 54.455 696.610 54.835 ;
        RECT 698.015 54.455 698.395 54.835 ;
        RECT 700.870 54.455 701.250 54.835 ;
        RECT 702.655 54.455 703.035 54.835 ;
        RECT 705.510 54.455 705.890 54.835 ;
        RECT 707.295 54.455 707.675 54.835 ;
        RECT 710.150 54.455 710.530 54.835 ;
        RECT 711.935 54.455 712.315 54.835 ;
        RECT 714.790 54.455 715.170 54.835 ;
        RECT 716.575 54.455 716.955 54.835 ;
        RECT 680.465 53.465 680.845 53.845 ;
        RECT 682.310 53.795 682.690 54.175 ;
        RECT 684.095 53.795 684.475 54.175 ;
        RECT 686.950 53.795 687.330 54.175 ;
        RECT 688.735 53.795 689.115 54.175 ;
        RECT 691.590 53.795 691.970 54.175 ;
        RECT 693.375 53.795 693.755 54.175 ;
        RECT 696.230 53.795 696.610 54.175 ;
        RECT 698.015 53.795 698.395 54.175 ;
        RECT 700.870 53.795 701.250 54.175 ;
        RECT 702.655 53.795 703.035 54.175 ;
        RECT 705.510 53.795 705.890 54.175 ;
        RECT 707.295 53.795 707.675 54.175 ;
        RECT 710.150 53.795 710.530 54.175 ;
        RECT 711.935 53.795 712.315 54.175 ;
        RECT 714.790 53.795 715.170 54.175 ;
        RECT 716.575 53.795 716.955 54.175 ;
        RECT 680.465 52.805 680.845 53.185 ;
        RECT 682.310 53.135 682.690 53.515 ;
        RECT 684.095 53.135 684.475 53.515 ;
        RECT 686.950 53.135 687.330 53.515 ;
        RECT 688.735 53.135 689.115 53.515 ;
        RECT 691.590 53.135 691.970 53.515 ;
        RECT 693.375 53.135 693.755 53.515 ;
        RECT 696.230 53.135 696.610 53.515 ;
        RECT 698.015 53.135 698.395 53.515 ;
        RECT 700.870 53.135 701.250 53.515 ;
        RECT 702.655 53.135 703.035 53.515 ;
        RECT 705.510 53.135 705.890 53.515 ;
        RECT 707.295 53.135 707.675 53.515 ;
        RECT 710.150 53.135 710.530 53.515 ;
        RECT 711.935 53.135 712.315 53.515 ;
        RECT 714.790 53.135 715.170 53.515 ;
        RECT 716.575 53.135 716.955 53.515 ;
        RECT 680.465 52.145 680.845 52.525 ;
        RECT 682.310 52.475 682.690 52.855 ;
        RECT 684.095 52.475 684.475 52.855 ;
        RECT 686.950 52.475 687.330 52.855 ;
        RECT 688.735 52.475 689.115 52.855 ;
        RECT 691.590 52.475 691.970 52.855 ;
        RECT 693.375 52.475 693.755 52.855 ;
        RECT 696.230 52.475 696.610 52.855 ;
        RECT 698.015 52.475 698.395 52.855 ;
        RECT 700.870 52.475 701.250 52.855 ;
        RECT 702.655 52.475 703.035 52.855 ;
        RECT 705.510 52.475 705.890 52.855 ;
        RECT 707.295 52.475 707.675 52.855 ;
        RECT 710.150 52.475 710.530 52.855 ;
        RECT 711.935 52.475 712.315 52.855 ;
        RECT 714.790 52.475 715.170 52.855 ;
        RECT 716.575 52.475 716.955 52.855 ;
        RECT 680.465 51.485 680.845 51.865 ;
        RECT 682.310 51.815 682.690 52.195 ;
        RECT 684.095 51.815 684.475 52.195 ;
        RECT 686.950 51.815 687.330 52.195 ;
        RECT 688.735 51.815 689.115 52.195 ;
        RECT 691.590 51.815 691.970 52.195 ;
        RECT 693.375 51.815 693.755 52.195 ;
        RECT 696.230 51.815 696.610 52.195 ;
        RECT 698.015 51.815 698.395 52.195 ;
        RECT 700.870 51.815 701.250 52.195 ;
        RECT 702.655 51.815 703.035 52.195 ;
        RECT 705.510 51.815 705.890 52.195 ;
        RECT 707.295 51.815 707.675 52.195 ;
        RECT 710.150 51.815 710.530 52.195 ;
        RECT 711.935 51.815 712.315 52.195 ;
        RECT 714.790 51.815 715.170 52.195 ;
        RECT 716.575 51.815 716.955 52.195 ;
        RECT 680.465 50.825 680.845 51.205 ;
        RECT 682.310 51.155 682.690 51.535 ;
        RECT 684.095 51.155 684.475 51.535 ;
        RECT 686.950 51.155 687.330 51.535 ;
        RECT 688.735 51.155 689.115 51.535 ;
        RECT 691.590 51.155 691.970 51.535 ;
        RECT 693.375 51.155 693.755 51.535 ;
        RECT 696.230 51.155 696.610 51.535 ;
        RECT 698.015 51.155 698.395 51.535 ;
        RECT 700.870 51.155 701.250 51.535 ;
        RECT 702.655 51.155 703.035 51.535 ;
        RECT 705.510 51.155 705.890 51.535 ;
        RECT 707.295 51.155 707.675 51.535 ;
        RECT 710.150 51.155 710.530 51.535 ;
        RECT 711.935 51.155 712.315 51.535 ;
        RECT 714.790 51.155 715.170 51.535 ;
        RECT 716.575 51.155 716.955 51.535 ;
        RECT 680.465 50.165 680.845 50.545 ;
        RECT 682.310 50.495 682.690 50.875 ;
        RECT 684.095 50.495 684.475 50.875 ;
        RECT 686.950 50.495 687.330 50.875 ;
        RECT 688.735 50.495 689.115 50.875 ;
        RECT 691.590 50.495 691.970 50.875 ;
        RECT 693.375 50.495 693.755 50.875 ;
        RECT 696.230 50.495 696.610 50.875 ;
        RECT 698.015 50.495 698.395 50.875 ;
        RECT 700.870 50.495 701.250 50.875 ;
        RECT 702.655 50.495 703.035 50.875 ;
        RECT 705.510 50.495 705.890 50.875 ;
        RECT 707.295 50.495 707.675 50.875 ;
        RECT 710.150 50.495 710.530 50.875 ;
        RECT 711.935 50.495 712.315 50.875 ;
        RECT 714.790 50.495 715.170 50.875 ;
        RECT 716.575 50.495 716.955 50.875 ;
        RECT 683.070 47.805 683.450 48.185 ;
        RECT 683.070 47.145 683.450 47.525 ;
        RECT 683.070 46.485 683.450 46.865 ;
        RECT 696.990 45.105 697.370 45.485 ;
        RECT 696.990 44.445 697.370 44.825 ;
        RECT 696.990 43.785 697.370 44.165 ;
        RECT 701.630 42.405 702.010 42.785 ;
        RECT 701.630 41.745 702.010 42.125 ;
        RECT 701.630 41.085 702.010 41.465 ;
        RECT 674.675 39.705 675.055 40.085 ;
        RECT 675.335 39.705 675.715 40.085 ;
        RECT 675.995 39.705 676.375 40.085 ;
        RECT 715.550 39.705 715.930 40.085 ;
        RECT 674.675 39.045 675.055 39.425 ;
        RECT 675.335 39.045 675.715 39.425 ;
        RECT 675.995 39.045 676.375 39.425 ;
        RECT 715.550 39.045 715.930 39.425 ;
        RECT 674.675 38.385 675.055 38.765 ;
        RECT 675.335 38.385 675.715 38.765 ;
        RECT 675.995 38.385 676.375 38.765 ;
        RECT 715.550 38.385 715.930 38.765 ;
        RECT 674.675 30.305 675.055 30.685 ;
        RECT 675.335 30.305 675.715 30.685 ;
        RECT 675.995 30.305 676.375 30.685 ;
        RECT 710.910 30.305 711.290 30.685 ;
        RECT 674.675 29.645 675.055 30.025 ;
        RECT 675.335 29.645 675.715 30.025 ;
        RECT 675.995 29.645 676.375 30.025 ;
        RECT 710.910 29.645 711.290 30.025 ;
        RECT 674.675 28.985 675.055 29.365 ;
        RECT 675.335 28.985 675.715 29.365 ;
        RECT 675.995 28.985 676.375 29.365 ;
        RECT 710.910 28.985 711.290 29.365 ;
        RECT 706.270 27.605 706.650 27.985 ;
        RECT 706.270 26.945 706.650 27.325 ;
        RECT 706.270 26.285 706.650 26.665 ;
        RECT 692.350 24.905 692.730 25.285 ;
        RECT 692.350 24.245 692.730 24.625 ;
        RECT 692.350 23.585 692.730 23.965 ;
        RECT 687.710 22.205 688.090 22.585 ;
        RECT 687.710 21.545 688.090 21.925 ;
        RECT 687.710 20.885 688.090 21.265 ;
        RECT 682.310 18.115 682.690 18.495 ;
        RECT 684.095 18.115 684.475 18.495 ;
        RECT 686.950 18.115 687.330 18.495 ;
        RECT 688.735 18.115 689.115 18.495 ;
        RECT 691.590 18.115 691.970 18.495 ;
        RECT 693.375 18.115 693.755 18.495 ;
        RECT 696.230 18.115 696.610 18.495 ;
        RECT 698.015 18.115 698.395 18.495 ;
        RECT 700.870 18.115 701.250 18.495 ;
        RECT 702.655 18.115 703.035 18.495 ;
        RECT 705.510 18.115 705.890 18.495 ;
        RECT 707.295 18.115 707.675 18.495 ;
        RECT 710.150 18.115 710.530 18.495 ;
        RECT 711.935 18.115 712.315 18.495 ;
        RECT 714.790 18.115 715.170 18.495 ;
        RECT 716.575 18.115 716.955 18.495 ;
        RECT 682.310 17.455 682.690 17.835 ;
        RECT 684.095 17.455 684.475 17.835 ;
        RECT 686.950 17.455 687.330 17.835 ;
        RECT 688.735 17.455 689.115 17.835 ;
        RECT 691.590 17.455 691.970 17.835 ;
        RECT 693.375 17.455 693.755 17.835 ;
        RECT 696.230 17.455 696.610 17.835 ;
        RECT 698.015 17.455 698.395 17.835 ;
        RECT 700.870 17.455 701.250 17.835 ;
        RECT 702.655 17.455 703.035 17.835 ;
        RECT 705.510 17.455 705.890 17.835 ;
        RECT 707.295 17.455 707.675 17.835 ;
        RECT 710.150 17.455 710.530 17.835 ;
        RECT 711.935 17.455 712.315 17.835 ;
        RECT 714.790 17.455 715.170 17.835 ;
        RECT 716.575 17.455 716.955 17.835 ;
        RECT 682.310 16.795 682.690 17.175 ;
        RECT 684.095 16.795 684.475 17.175 ;
        RECT 686.950 16.795 687.330 17.175 ;
        RECT 688.735 16.795 689.115 17.175 ;
        RECT 691.590 16.795 691.970 17.175 ;
        RECT 693.375 16.795 693.755 17.175 ;
        RECT 696.230 16.795 696.610 17.175 ;
        RECT 698.015 16.795 698.395 17.175 ;
        RECT 700.870 16.795 701.250 17.175 ;
        RECT 702.655 16.795 703.035 17.175 ;
        RECT 705.510 16.795 705.890 17.175 ;
        RECT 707.295 16.795 707.675 17.175 ;
        RECT 710.150 16.795 710.530 17.175 ;
        RECT 711.935 16.795 712.315 17.175 ;
        RECT 714.790 16.795 715.170 17.175 ;
        RECT 716.575 16.795 716.955 17.175 ;
        RECT 682.310 16.135 682.690 16.515 ;
        RECT 684.095 16.135 684.475 16.515 ;
        RECT 686.950 16.135 687.330 16.515 ;
        RECT 688.735 16.135 689.115 16.515 ;
        RECT 691.590 16.135 691.970 16.515 ;
        RECT 693.375 16.135 693.755 16.515 ;
        RECT 696.230 16.135 696.610 16.515 ;
        RECT 698.015 16.135 698.395 16.515 ;
        RECT 700.870 16.135 701.250 16.515 ;
        RECT 702.655 16.135 703.035 16.515 ;
        RECT 705.510 16.135 705.890 16.515 ;
        RECT 707.295 16.135 707.675 16.515 ;
        RECT 710.150 16.135 710.530 16.515 ;
        RECT 711.935 16.135 712.315 16.515 ;
        RECT 714.790 16.135 715.170 16.515 ;
        RECT 716.575 16.135 716.955 16.515 ;
        RECT 682.310 15.475 682.690 15.855 ;
        RECT 684.095 15.475 684.475 15.855 ;
        RECT 686.950 15.475 687.330 15.855 ;
        RECT 688.735 15.475 689.115 15.855 ;
        RECT 691.590 15.475 691.970 15.855 ;
        RECT 693.375 15.475 693.755 15.855 ;
        RECT 696.230 15.475 696.610 15.855 ;
        RECT 698.015 15.475 698.395 15.855 ;
        RECT 700.870 15.475 701.250 15.855 ;
        RECT 702.655 15.475 703.035 15.855 ;
        RECT 705.510 15.475 705.890 15.855 ;
        RECT 707.295 15.475 707.675 15.855 ;
        RECT 710.150 15.475 710.530 15.855 ;
        RECT 711.935 15.475 712.315 15.855 ;
        RECT 714.790 15.475 715.170 15.855 ;
        RECT 716.575 15.475 716.955 15.855 ;
        RECT 682.310 14.815 682.690 15.195 ;
        RECT 684.095 14.815 684.475 15.195 ;
        RECT 686.950 14.815 687.330 15.195 ;
        RECT 688.735 14.815 689.115 15.195 ;
        RECT 691.590 14.815 691.970 15.195 ;
        RECT 693.375 14.815 693.755 15.195 ;
        RECT 696.230 14.815 696.610 15.195 ;
        RECT 698.015 14.815 698.395 15.195 ;
        RECT 700.870 14.815 701.250 15.195 ;
        RECT 702.655 14.815 703.035 15.195 ;
        RECT 705.510 14.815 705.890 15.195 ;
        RECT 707.295 14.815 707.675 15.195 ;
        RECT 710.150 14.815 710.530 15.195 ;
        RECT 711.935 14.815 712.315 15.195 ;
        RECT 714.790 14.815 715.170 15.195 ;
        RECT 716.575 14.815 716.955 15.195 ;
        RECT 682.310 14.155 682.690 14.535 ;
        RECT 684.095 14.155 684.475 14.535 ;
        RECT 686.950 14.155 687.330 14.535 ;
        RECT 688.735 14.155 689.115 14.535 ;
        RECT 691.590 14.155 691.970 14.535 ;
        RECT 693.375 14.155 693.755 14.535 ;
        RECT 696.230 14.155 696.610 14.535 ;
        RECT 698.015 14.155 698.395 14.535 ;
        RECT 700.870 14.155 701.250 14.535 ;
        RECT 702.655 14.155 703.035 14.535 ;
        RECT 705.510 14.155 705.890 14.535 ;
        RECT 707.295 14.155 707.675 14.535 ;
        RECT 710.150 14.155 710.530 14.535 ;
        RECT 711.935 14.155 712.315 14.535 ;
        RECT 714.790 14.155 715.170 14.535 ;
        RECT 716.575 14.155 716.955 14.535 ;
        RECT 682.310 13.495 682.690 13.875 ;
        RECT 684.095 13.495 684.475 13.875 ;
        RECT 686.950 13.495 687.330 13.875 ;
        RECT 688.735 13.495 689.115 13.875 ;
        RECT 691.590 13.495 691.970 13.875 ;
        RECT 693.375 13.495 693.755 13.875 ;
        RECT 696.230 13.495 696.610 13.875 ;
        RECT 698.015 13.495 698.395 13.875 ;
        RECT 700.870 13.495 701.250 13.875 ;
        RECT 702.655 13.495 703.035 13.875 ;
        RECT 705.510 13.495 705.890 13.875 ;
        RECT 707.295 13.495 707.675 13.875 ;
        RECT 710.150 13.495 710.530 13.875 ;
        RECT 711.935 13.495 712.315 13.875 ;
        RECT 714.790 13.495 715.170 13.875 ;
        RECT 716.575 13.495 716.955 13.875 ;
        RECT 682.310 12.835 682.690 13.215 ;
        RECT 684.095 12.835 684.475 13.215 ;
        RECT 686.950 12.835 687.330 13.215 ;
        RECT 688.735 12.835 689.115 13.215 ;
        RECT 691.590 12.835 691.970 13.215 ;
        RECT 693.375 12.835 693.755 13.215 ;
        RECT 696.230 12.835 696.610 13.215 ;
        RECT 698.015 12.835 698.395 13.215 ;
        RECT 700.870 12.835 701.250 13.215 ;
        RECT 702.655 12.835 703.035 13.215 ;
        RECT 705.510 12.835 705.890 13.215 ;
        RECT 707.295 12.835 707.675 13.215 ;
        RECT 710.150 12.835 710.530 13.215 ;
        RECT 711.935 12.835 712.315 13.215 ;
        RECT 714.790 12.835 715.170 13.215 ;
        RECT 716.575 12.835 716.955 13.215 ;
        RECT 682.310 12.175 682.690 12.555 ;
        RECT 684.095 12.175 684.475 12.555 ;
        RECT 686.950 12.175 687.330 12.555 ;
        RECT 688.735 12.175 689.115 12.555 ;
        RECT 691.590 12.175 691.970 12.555 ;
        RECT 693.375 12.175 693.755 12.555 ;
        RECT 696.230 12.175 696.610 12.555 ;
        RECT 698.015 12.175 698.395 12.555 ;
        RECT 700.870 12.175 701.250 12.555 ;
        RECT 702.655 12.175 703.035 12.555 ;
        RECT 705.510 12.175 705.890 12.555 ;
        RECT 707.295 12.175 707.675 12.555 ;
        RECT 710.150 12.175 710.530 12.555 ;
        RECT 711.935 12.175 712.315 12.555 ;
        RECT 714.790 12.175 715.170 12.555 ;
        RECT 716.575 12.175 716.955 12.555 ;
        RECT 682.310 11.515 682.690 11.895 ;
        RECT 684.095 11.515 684.475 11.895 ;
        RECT 686.950 11.515 687.330 11.895 ;
        RECT 688.735 11.515 689.115 11.895 ;
        RECT 691.590 11.515 691.970 11.895 ;
        RECT 693.375 11.515 693.755 11.895 ;
        RECT 696.230 11.515 696.610 11.895 ;
        RECT 698.015 11.515 698.395 11.895 ;
        RECT 700.870 11.515 701.250 11.895 ;
        RECT 702.655 11.515 703.035 11.895 ;
        RECT 705.510 11.515 705.890 11.895 ;
        RECT 707.295 11.515 707.675 11.895 ;
        RECT 710.150 11.515 710.530 11.895 ;
        RECT 711.935 11.515 712.315 11.895 ;
        RECT 714.790 11.515 715.170 11.895 ;
        RECT 716.575 11.515 716.955 11.895 ;
        RECT 682.310 10.855 682.690 11.235 ;
        RECT 684.095 10.855 684.475 11.235 ;
        RECT 686.950 10.855 687.330 11.235 ;
        RECT 688.735 10.855 689.115 11.235 ;
        RECT 691.590 10.855 691.970 11.235 ;
        RECT 693.375 10.855 693.755 11.235 ;
        RECT 696.230 10.855 696.610 11.235 ;
        RECT 698.015 10.855 698.395 11.235 ;
        RECT 700.870 10.855 701.250 11.235 ;
        RECT 702.655 10.855 703.035 11.235 ;
        RECT 705.510 10.855 705.890 11.235 ;
        RECT 707.295 10.855 707.675 11.235 ;
        RECT 710.150 10.855 710.530 11.235 ;
        RECT 711.935 10.855 712.315 11.235 ;
        RECT 714.790 10.855 715.170 11.235 ;
        RECT 716.575 10.855 716.955 11.235 ;
        RECT 682.310 10.195 682.690 10.575 ;
        RECT 684.095 10.195 684.475 10.575 ;
        RECT 686.950 10.195 687.330 10.575 ;
        RECT 688.735 10.195 689.115 10.575 ;
        RECT 691.590 10.195 691.970 10.575 ;
        RECT 693.375 10.195 693.755 10.575 ;
        RECT 696.230 10.195 696.610 10.575 ;
        RECT 698.015 10.195 698.395 10.575 ;
        RECT 700.870 10.195 701.250 10.575 ;
        RECT 702.655 10.195 703.035 10.575 ;
        RECT 705.510 10.195 705.890 10.575 ;
        RECT 707.295 10.195 707.675 10.575 ;
        RECT 710.150 10.195 710.530 10.575 ;
        RECT 711.935 10.195 712.315 10.575 ;
        RECT 714.790 10.195 715.170 10.575 ;
        RECT 716.575 10.195 716.955 10.575 ;
        RECT 682.310 9.535 682.690 9.915 ;
        RECT 684.095 9.535 684.475 9.915 ;
        RECT 686.950 9.535 687.330 9.915 ;
        RECT 688.735 9.535 689.115 9.915 ;
        RECT 691.590 9.535 691.970 9.915 ;
        RECT 693.375 9.535 693.755 9.915 ;
        RECT 696.230 9.535 696.610 9.915 ;
        RECT 698.015 9.535 698.395 9.915 ;
        RECT 700.870 9.535 701.250 9.915 ;
        RECT 702.655 9.535 703.035 9.915 ;
        RECT 705.510 9.535 705.890 9.915 ;
        RECT 707.295 9.535 707.675 9.915 ;
        RECT 710.150 9.535 710.530 9.915 ;
        RECT 711.935 9.535 712.315 9.915 ;
        RECT 714.790 9.535 715.170 9.915 ;
        RECT 716.575 9.535 716.955 9.915 ;
        RECT 647.550 8.770 653.955 9.100 ;
        RECT 647.550 8.750 651.515 8.770 ;
        RECT 611.190 4.690 611.570 5.070 ;
        RECT 612.190 4.690 612.570 5.070 ;
        RECT 612.850 4.690 613.230 5.070 ;
        RECT 613.510 4.690 613.890 5.070 ;
        RECT 614.430 4.690 614.810 5.070 ;
        RECT 615.090 4.690 615.470 5.070 ;
        RECT 615.750 4.690 616.130 5.070 ;
        RECT 616.670 4.690 617.050 5.070 ;
        RECT 617.330 4.690 617.710 5.070 ;
        RECT 617.990 4.690 618.370 5.070 ;
        RECT 618.910 4.690 619.290 5.070 ;
        RECT 619.570 4.690 619.950 5.070 ;
        RECT 620.230 4.690 620.610 5.070 ;
        RECT 621.150 4.690 621.530 5.070 ;
        RECT 621.810 4.690 622.190 5.070 ;
        RECT 622.470 4.690 622.850 5.070 ;
        RECT 623.390 4.690 623.770 5.070 ;
        RECT 624.050 4.690 624.430 5.070 ;
        RECT 624.710 4.690 625.090 5.070 ;
        RECT 625.630 4.690 626.010 5.070 ;
        RECT 626.290 4.690 626.670 5.070 ;
        RECT 626.950 4.690 627.330 5.070 ;
        RECT 627.870 4.690 628.250 5.070 ;
        RECT 628.530 4.690 628.910 5.070 ;
        RECT 629.190 4.690 629.570 5.070 ;
        RECT 630.110 4.690 630.490 5.070 ;
        RECT 630.770 4.690 631.150 5.070 ;
        RECT 631.430 4.690 631.810 5.070 ;
        RECT 632.470 4.690 632.850 5.070 ;
        RECT 633.470 4.690 633.850 5.070 ;
        RECT 634.130 4.690 634.510 5.070 ;
        RECT 634.790 4.690 635.170 5.070 ;
        RECT 635.710 4.690 636.090 5.070 ;
        RECT 636.370 4.690 636.750 5.070 ;
        RECT 637.030 4.690 637.410 5.070 ;
        RECT 637.950 4.690 638.330 5.070 ;
        RECT 638.610 4.690 638.990 5.070 ;
        RECT 639.270 4.690 639.650 5.070 ;
        RECT 640.190 4.690 640.570 5.070 ;
        RECT 640.850 4.690 641.230 5.070 ;
        RECT 641.510 4.690 641.890 5.070 ;
        RECT 642.430 4.690 642.810 5.070 ;
        RECT 643.090 4.690 643.470 5.070 ;
        RECT 643.750 4.690 644.130 5.070 ;
        RECT 644.670 4.690 645.050 5.070 ;
        RECT 645.330 4.690 645.710 5.070 ;
        RECT 645.990 4.690 646.370 5.070 ;
        RECT 646.910 4.690 647.290 5.070 ;
        RECT 647.570 4.690 647.950 5.070 ;
        RECT 648.230 4.690 648.610 5.070 ;
        RECT 649.150 4.690 649.530 5.070 ;
        RECT 649.810 4.690 650.190 5.070 ;
        RECT 650.470 4.690 650.850 5.070 ;
        RECT 651.490 4.690 651.870 5.070 ;
        RECT 652.150 4.690 652.530 5.070 ;
        RECT 652.810 4.690 653.190 5.070 ;
        RECT 653.625 4.150 653.955 8.770 ;
        RECT 668.125 8.750 672.090 9.150 ;
        RECT 682.310 8.875 682.690 9.255 ;
        RECT 684.095 8.875 684.475 9.255 ;
        RECT 686.950 8.875 687.330 9.255 ;
        RECT 688.735 8.875 689.115 9.255 ;
        RECT 691.590 8.875 691.970 9.255 ;
        RECT 693.375 8.875 693.755 9.255 ;
        RECT 696.230 8.875 696.610 9.255 ;
        RECT 698.015 8.875 698.395 9.255 ;
        RECT 700.870 8.875 701.250 9.255 ;
        RECT 702.655 8.875 703.035 9.255 ;
        RECT 705.510 8.875 705.890 9.255 ;
        RECT 707.295 8.875 707.675 9.255 ;
        RECT 710.150 8.875 710.530 9.255 ;
        RECT 711.935 8.875 712.315 9.255 ;
        RECT 714.790 8.875 715.170 9.255 ;
        RECT 716.575 8.875 716.955 9.255 ;
        RECT 654.870 4.690 655.250 5.070 ;
        RECT 655.870 4.690 656.250 5.070 ;
        RECT 656.530 4.690 656.910 5.070 ;
        RECT 657.190 4.690 657.570 5.070 ;
        RECT 658.110 4.690 658.490 5.070 ;
        RECT 658.770 4.690 659.150 5.070 ;
        RECT 659.430 4.690 659.810 5.070 ;
        RECT 660.350 4.690 660.730 5.070 ;
        RECT 661.010 4.690 661.390 5.070 ;
        RECT 661.670 4.690 662.050 5.070 ;
        RECT 662.590 4.690 662.970 5.070 ;
        RECT 663.250 4.690 663.630 5.070 ;
        RECT 663.910 4.690 664.290 5.070 ;
        RECT 664.830 4.690 665.210 5.070 ;
        RECT 665.490 4.690 665.870 5.070 ;
        RECT 666.150 4.690 666.530 5.070 ;
        RECT 667.070 4.690 667.450 5.070 ;
        RECT 667.730 4.690 668.110 5.070 ;
        RECT 668.390 4.690 668.770 5.070 ;
        RECT 669.310 4.690 669.690 5.070 ;
        RECT 669.970 4.690 670.350 5.070 ;
        RECT 670.630 4.690 671.010 5.070 ;
        RECT 671.550 4.690 671.930 5.070 ;
        RECT 672.210 4.690 672.590 5.070 ;
        RECT 672.870 4.690 673.250 5.070 ;
        RECT 673.790 4.690 674.170 5.070 ;
        RECT 674.450 4.690 674.830 5.070 ;
        RECT 675.110 4.690 675.490 5.070 ;
        RECT 676.150 4.690 676.530 5.070 ;
        RECT 677.150 4.690 677.530 5.070 ;
        RECT 677.810 4.690 678.190 5.070 ;
        RECT 678.470 4.690 678.850 5.070 ;
        RECT 679.490 4.690 679.870 5.070 ;
        RECT 121.420 3.420 121.800 3.800 ;
        RECT 142.880 3.770 143.260 4.150 ;
        RECT 184.320 3.770 184.700 4.150 ;
        RECT 228.000 3.770 228.380 4.150 ;
        RECT 269.440 3.770 269.820 4.150 ;
        RECT 313.120 3.770 313.500 4.150 ;
        RECT 354.560 3.770 354.940 4.150 ;
        RECT 398.240 3.770 398.620 4.150 ;
        RECT 439.680 3.770 440.060 4.150 ;
        RECT 483.360 3.770 483.740 4.150 ;
        RECT 524.800 3.770 525.180 4.150 ;
        RECT 568.480 3.770 568.860 4.150 ;
        RECT 609.920 3.770 610.300 4.150 ;
        RECT 653.600 3.770 653.980 4.150 ;
        RECT 120.740 2.580 121.440 2.950 ;
        RECT 121.830 2.760 122.210 3.140 ;
        RECT 124.245 2.950 127.455 3.300 ;
        RECT 121.070 2.305 121.440 2.580 ;
        RECT 124.245 2.305 124.595 2.950 ;
        RECT 128.730 2.760 130.250 3.255 ;
        RECT 132.195 3.125 132.575 3.150 ;
        RECT 131.115 2.795 132.575 3.125 ;
        RECT 128.730 2.600 129.140 2.760 ;
        RECT 121.070 1.955 124.595 2.305 ;
        RECT 124.895 2.250 129.140 2.600 ;
        RECT 114.510 1.555 116.615 1.885 ;
        RECT 129.340 1.885 129.720 1.910 ;
        RECT 131.115 1.885 131.445 2.795 ;
        RECT 132.195 2.770 132.575 2.795 ;
        RECT 129.340 1.555 131.445 1.885 ;
        RECT 12.090 1.530 12.470 1.555 ;
        RECT 30.280 1.530 30.660 1.555 ;
        RECT 46.230 1.530 46.610 1.555 ;
        RECT 61.060 1.530 61.440 1.555 ;
        RECT 80.370 1.530 80.750 1.555 ;
        RECT 95.200 1.530 95.580 1.555 ;
        RECT 114.510 1.530 114.890 1.555 ;
        RECT 129.340 1.530 129.720 1.555 ;
        RECT 0.850 0.770 1.230 1.150 ;
        RECT 1.990 0.770 2.370 1.150 ;
        RECT 7.430 0.770 7.810 1.150 ;
        RECT 8.090 0.770 8.470 1.150 ;
        RECT 8.750 0.770 9.130 1.150 ;
        RECT 14.300 0.770 14.680 1.150 ;
        RECT 15.620 0.770 16.000 1.150 ;
        RECT 17.660 0.770 18.040 1.150 ;
        RECT 18.980 0.770 19.360 1.150 ;
        RECT 25.620 0.770 26.000 1.150 ;
        RECT 26.280 0.770 26.660 1.150 ;
        RECT 26.940 0.770 27.320 1.150 ;
        RECT 32.490 0.770 32.870 1.150 ;
        RECT 33.810 0.770 34.190 1.150 ;
        RECT 36.130 0.770 36.510 1.150 ;
        RECT 41.570 0.770 41.950 1.150 ;
        RECT 42.230 0.770 42.610 1.150 ;
        RECT 42.890 0.770 43.270 1.150 ;
        RECT 48.440 0.770 48.820 1.150 ;
        RECT 49.760 0.770 50.140 1.150 ;
        RECT 56.400 0.770 56.780 1.150 ;
        RECT 57.060 0.770 57.440 1.150 ;
        RECT 57.720 0.770 58.100 1.150 ;
        RECT 63.270 0.770 63.650 1.150 ;
        RECT 64.590 0.770 64.970 1.150 ;
        RECT 66.630 0.770 67.010 1.150 ;
        RECT 67.950 0.770 68.330 1.150 ;
        RECT 70.270 0.770 70.650 1.150 ;
        RECT 75.710 0.770 76.090 1.150 ;
        RECT 76.370 0.770 76.750 1.150 ;
        RECT 77.030 0.770 77.410 1.150 ;
        RECT 82.580 0.770 82.960 1.150 ;
        RECT 83.900 0.770 84.280 1.150 ;
        RECT 90.540 0.770 90.920 1.150 ;
        RECT 91.200 0.770 91.580 1.150 ;
        RECT 91.860 0.770 92.240 1.150 ;
        RECT 97.410 0.770 97.790 1.150 ;
        RECT 98.730 0.770 99.110 1.150 ;
        RECT 100.770 0.770 101.150 1.150 ;
        RECT 102.090 0.770 102.470 1.150 ;
        RECT 104.410 0.770 104.790 1.150 ;
        RECT 109.850 0.770 110.230 1.150 ;
        RECT 110.510 0.770 110.890 1.150 ;
        RECT 111.170 0.770 111.550 1.150 ;
        RECT 116.720 0.770 117.100 1.150 ;
        RECT 118.040 0.770 118.420 1.150 ;
        RECT 124.680 0.770 125.060 1.150 ;
        RECT 125.340 0.770 125.720 1.150 ;
        RECT 126.000 0.770 126.380 1.150 ;
        RECT 131.550 0.770 131.930 1.150 ;
        RECT 132.870 0.770 133.250 1.150 ;
        RECT 135.190 0.770 135.570 1.150 ;
        RECT 136.190 0.770 136.570 1.150 ;
        RECT 136.850 0.770 137.230 1.150 ;
        RECT 137.510 0.770 137.890 1.150 ;
        RECT 138.430 0.770 138.810 1.150 ;
        RECT 139.090 0.770 139.470 1.150 ;
        RECT 139.750 0.770 140.130 1.150 ;
        RECT 140.510 0.770 140.890 1.150 ;
        RECT 141.830 0.770 142.210 1.150 ;
        RECT 144.030 0.770 144.410 1.150 ;
        RECT 144.690 0.770 145.070 1.150 ;
        RECT 145.350 0.770 145.730 1.150 ;
        RECT 146.270 0.770 146.650 1.150 ;
        RECT 146.930 0.770 147.310 1.150 ;
        RECT 147.590 0.770 147.970 1.150 ;
        RECT 148.510 0.770 148.890 1.150 ;
        RECT 149.170 0.770 149.550 1.150 ;
        RECT 149.830 0.770 150.210 1.150 ;
        RECT 150.750 0.770 151.130 1.150 ;
        RECT 151.410 0.770 151.790 1.150 ;
        RECT 152.070 0.770 152.450 1.150 ;
        RECT 152.990 0.770 153.370 1.150 ;
        RECT 153.650 0.770 154.030 1.150 ;
        RECT 154.310 0.770 154.690 1.150 ;
        RECT 155.350 0.770 155.730 1.150 ;
        RECT 156.350 0.770 156.730 1.150 ;
        RECT 157.010 0.770 157.390 1.150 ;
        RECT 157.670 0.770 158.050 1.150 ;
        RECT 158.590 0.770 158.970 1.150 ;
        RECT 159.250 0.770 159.630 1.150 ;
        RECT 159.910 0.770 160.290 1.150 ;
        RECT 160.830 0.770 161.210 1.150 ;
        RECT 161.490 0.770 161.870 1.150 ;
        RECT 162.150 0.770 162.530 1.150 ;
        RECT 163.070 0.770 163.450 1.150 ;
        RECT 163.730 0.770 164.110 1.150 ;
        RECT 164.390 0.770 164.770 1.150 ;
        RECT 165.310 0.770 165.690 1.150 ;
        RECT 165.970 0.770 166.350 1.150 ;
        RECT 166.630 0.770 167.010 1.150 ;
        RECT 167.550 0.770 167.930 1.150 ;
        RECT 168.210 0.770 168.590 1.150 ;
        RECT 168.870 0.770 169.250 1.150 ;
        RECT 169.790 0.770 170.170 1.150 ;
        RECT 170.450 0.770 170.830 1.150 ;
        RECT 171.110 0.770 171.490 1.150 ;
        RECT 172.030 0.770 172.410 1.150 ;
        RECT 172.690 0.770 173.070 1.150 ;
        RECT 173.350 0.770 173.730 1.150 ;
        RECT 174.270 0.770 174.650 1.150 ;
        RECT 174.930 0.770 175.310 1.150 ;
        RECT 175.590 0.770 175.970 1.150 ;
        RECT 176.630 0.770 177.010 1.150 ;
        RECT 177.630 0.770 178.010 1.150 ;
        RECT 178.290 0.770 178.670 1.150 ;
        RECT 178.950 0.770 179.330 1.150 ;
        RECT 179.870 0.770 180.250 1.150 ;
        RECT 180.530 0.770 180.910 1.150 ;
        RECT 181.190 0.770 181.570 1.150 ;
        RECT 181.950 0.770 182.330 1.150 ;
        RECT 183.270 0.770 183.650 1.150 ;
        RECT 185.470 0.770 185.850 1.150 ;
        RECT 186.130 0.770 186.510 1.150 ;
        RECT 186.790 0.770 187.170 1.150 ;
        RECT 187.710 0.770 188.090 1.150 ;
        RECT 188.370 0.770 188.750 1.150 ;
        RECT 189.030 0.770 189.410 1.150 ;
        RECT 189.950 0.770 190.330 1.150 ;
        RECT 190.610 0.770 190.990 1.150 ;
        RECT 191.270 0.770 191.650 1.150 ;
        RECT 192.190 0.770 192.570 1.150 ;
        RECT 192.850 0.770 193.230 1.150 ;
        RECT 193.510 0.770 193.890 1.150 ;
        RECT 194.430 0.770 194.810 1.150 ;
        RECT 195.090 0.770 195.470 1.150 ;
        RECT 195.750 0.770 196.130 1.150 ;
        RECT 196.790 0.770 197.170 1.150 ;
        RECT 197.790 0.770 198.170 1.150 ;
        RECT 198.450 0.770 198.830 1.150 ;
        RECT 199.110 0.770 199.490 1.150 ;
        RECT 200.030 0.770 200.410 1.150 ;
        RECT 200.690 0.770 201.070 1.150 ;
        RECT 201.350 0.770 201.730 1.150 ;
        RECT 202.270 0.770 202.650 1.150 ;
        RECT 202.930 0.770 203.310 1.150 ;
        RECT 203.590 0.770 203.970 1.150 ;
        RECT 204.510 0.770 204.890 1.150 ;
        RECT 205.170 0.770 205.550 1.150 ;
        RECT 205.830 0.770 206.210 1.150 ;
        RECT 206.750 0.770 207.130 1.150 ;
        RECT 207.410 0.770 207.790 1.150 ;
        RECT 208.070 0.770 208.450 1.150 ;
        RECT 208.990 0.770 209.370 1.150 ;
        RECT 209.650 0.770 210.030 1.150 ;
        RECT 210.310 0.770 210.690 1.150 ;
        RECT 211.230 0.770 211.610 1.150 ;
        RECT 211.890 0.770 212.270 1.150 ;
        RECT 212.550 0.770 212.930 1.150 ;
        RECT 213.470 0.770 213.850 1.150 ;
        RECT 214.130 0.770 214.510 1.150 ;
        RECT 214.790 0.770 215.170 1.150 ;
        RECT 215.710 0.770 216.090 1.150 ;
        RECT 216.370 0.770 216.750 1.150 ;
        RECT 217.030 0.770 217.410 1.150 ;
        RECT 218.070 0.770 218.450 1.150 ;
        RECT 219.070 0.770 219.450 1.150 ;
        RECT 219.730 0.770 220.110 1.150 ;
        RECT 220.390 0.770 220.770 1.150 ;
        RECT 221.310 0.770 221.690 1.150 ;
        RECT 221.970 0.770 222.350 1.150 ;
        RECT 222.630 0.770 223.010 1.150 ;
        RECT 223.550 0.770 223.930 1.150 ;
        RECT 224.210 0.770 224.590 1.150 ;
        RECT 224.870 0.770 225.250 1.150 ;
        RECT 225.630 0.770 226.010 1.150 ;
        RECT 226.950 0.770 227.330 1.150 ;
        RECT 229.150 0.770 229.530 1.150 ;
        RECT 229.810 0.770 230.190 1.150 ;
        RECT 230.470 0.770 230.850 1.150 ;
        RECT 231.390 0.770 231.770 1.150 ;
        RECT 232.050 0.770 232.430 1.150 ;
        RECT 232.710 0.770 233.090 1.150 ;
        RECT 233.630 0.770 234.010 1.150 ;
        RECT 234.290 0.770 234.670 1.150 ;
        RECT 234.950 0.770 235.330 1.150 ;
        RECT 235.870 0.770 236.250 1.150 ;
        RECT 236.530 0.770 236.910 1.150 ;
        RECT 237.190 0.770 237.570 1.150 ;
        RECT 238.230 0.770 238.610 1.150 ;
        RECT 239.230 0.770 239.610 1.150 ;
        RECT 239.890 0.770 240.270 1.150 ;
        RECT 240.550 0.770 240.930 1.150 ;
        RECT 241.470 0.770 241.850 1.150 ;
        RECT 242.130 0.770 242.510 1.150 ;
        RECT 242.790 0.770 243.170 1.150 ;
        RECT 243.710 0.770 244.090 1.150 ;
        RECT 244.370 0.770 244.750 1.150 ;
        RECT 245.030 0.770 245.410 1.150 ;
        RECT 245.950 0.770 246.330 1.150 ;
        RECT 246.610 0.770 246.990 1.150 ;
        RECT 247.270 0.770 247.650 1.150 ;
        RECT 248.190 0.770 248.570 1.150 ;
        RECT 248.850 0.770 249.230 1.150 ;
        RECT 249.510 0.770 249.890 1.150 ;
        RECT 250.430 0.770 250.810 1.150 ;
        RECT 251.090 0.770 251.470 1.150 ;
        RECT 251.750 0.770 252.130 1.150 ;
        RECT 252.670 0.770 253.050 1.150 ;
        RECT 253.330 0.770 253.710 1.150 ;
        RECT 253.990 0.770 254.370 1.150 ;
        RECT 254.910 0.770 255.290 1.150 ;
        RECT 255.570 0.770 255.950 1.150 ;
        RECT 256.230 0.770 256.610 1.150 ;
        RECT 257.150 0.770 257.530 1.150 ;
        RECT 257.810 0.770 258.190 1.150 ;
        RECT 258.470 0.770 258.850 1.150 ;
        RECT 259.510 0.770 259.890 1.150 ;
        RECT 260.510 0.770 260.890 1.150 ;
        RECT 261.170 0.770 261.550 1.150 ;
        RECT 261.830 0.770 262.210 1.150 ;
        RECT 262.750 0.770 263.130 1.150 ;
        RECT 263.410 0.770 263.790 1.150 ;
        RECT 264.070 0.770 264.450 1.150 ;
        RECT 264.990 0.770 265.370 1.150 ;
        RECT 265.650 0.770 266.030 1.150 ;
        RECT 266.310 0.770 266.690 1.150 ;
        RECT 267.070 0.770 267.450 1.150 ;
        RECT 268.390 0.770 268.770 1.150 ;
        RECT 270.590 0.770 270.970 1.150 ;
        RECT 271.250 0.770 271.630 1.150 ;
        RECT 271.910 0.770 272.290 1.150 ;
        RECT 272.830 0.770 273.210 1.150 ;
        RECT 273.490 0.770 273.870 1.150 ;
        RECT 274.150 0.770 274.530 1.150 ;
        RECT 275.070 0.770 275.450 1.150 ;
        RECT 275.730 0.770 276.110 1.150 ;
        RECT 276.390 0.770 276.770 1.150 ;
        RECT 277.310 0.770 277.690 1.150 ;
        RECT 277.970 0.770 278.350 1.150 ;
        RECT 278.630 0.770 279.010 1.150 ;
        RECT 279.670 0.770 280.050 1.150 ;
        RECT 280.670 0.770 281.050 1.150 ;
        RECT 281.330 0.770 281.710 1.150 ;
        RECT 281.990 0.770 282.370 1.150 ;
        RECT 282.910 0.770 283.290 1.150 ;
        RECT 283.570 0.770 283.950 1.150 ;
        RECT 284.230 0.770 284.610 1.150 ;
        RECT 285.150 0.770 285.530 1.150 ;
        RECT 285.810 0.770 286.190 1.150 ;
        RECT 286.470 0.770 286.850 1.150 ;
        RECT 287.390 0.770 287.770 1.150 ;
        RECT 288.050 0.770 288.430 1.150 ;
        RECT 288.710 0.770 289.090 1.150 ;
        RECT 289.630 0.770 290.010 1.150 ;
        RECT 290.290 0.770 290.670 1.150 ;
        RECT 290.950 0.770 291.330 1.150 ;
        RECT 291.870 0.770 292.250 1.150 ;
        RECT 292.530 0.770 292.910 1.150 ;
        RECT 293.190 0.770 293.570 1.150 ;
        RECT 294.110 0.770 294.490 1.150 ;
        RECT 294.770 0.770 295.150 1.150 ;
        RECT 295.430 0.770 295.810 1.150 ;
        RECT 296.350 0.770 296.730 1.150 ;
        RECT 297.010 0.770 297.390 1.150 ;
        RECT 297.670 0.770 298.050 1.150 ;
        RECT 298.590 0.770 298.970 1.150 ;
        RECT 299.250 0.770 299.630 1.150 ;
        RECT 299.910 0.770 300.290 1.150 ;
        RECT 300.950 0.770 301.330 1.150 ;
        RECT 301.950 0.770 302.330 1.150 ;
        RECT 302.610 0.770 302.990 1.150 ;
        RECT 303.270 0.770 303.650 1.150 ;
        RECT 304.190 0.770 304.570 1.150 ;
        RECT 304.850 0.770 305.230 1.150 ;
        RECT 305.510 0.770 305.890 1.150 ;
        RECT 306.430 0.770 306.810 1.150 ;
        RECT 307.090 0.770 307.470 1.150 ;
        RECT 307.750 0.770 308.130 1.150 ;
        RECT 308.670 0.770 309.050 1.150 ;
        RECT 309.330 0.770 309.710 1.150 ;
        RECT 309.990 0.770 310.370 1.150 ;
        RECT 310.750 0.770 311.130 1.150 ;
        RECT 312.070 0.770 312.450 1.150 ;
        RECT 314.270 0.770 314.650 1.150 ;
        RECT 314.930 0.770 315.310 1.150 ;
        RECT 315.590 0.770 315.970 1.150 ;
        RECT 316.510 0.770 316.890 1.150 ;
        RECT 317.170 0.770 317.550 1.150 ;
        RECT 317.830 0.770 318.210 1.150 ;
        RECT 318.750 0.770 319.130 1.150 ;
        RECT 319.410 0.770 319.790 1.150 ;
        RECT 320.070 0.770 320.450 1.150 ;
        RECT 321.110 0.770 321.490 1.150 ;
        RECT 322.110 0.770 322.490 1.150 ;
        RECT 322.770 0.770 323.150 1.150 ;
        RECT 323.430 0.770 323.810 1.150 ;
        RECT 324.350 0.770 324.730 1.150 ;
        RECT 325.010 0.770 325.390 1.150 ;
        RECT 325.670 0.770 326.050 1.150 ;
        RECT 326.590 0.770 326.970 1.150 ;
        RECT 327.250 0.770 327.630 1.150 ;
        RECT 327.910 0.770 328.290 1.150 ;
        RECT 328.830 0.770 329.210 1.150 ;
        RECT 329.490 0.770 329.870 1.150 ;
        RECT 330.150 0.770 330.530 1.150 ;
        RECT 331.070 0.770 331.450 1.150 ;
        RECT 331.730 0.770 332.110 1.150 ;
        RECT 332.390 0.770 332.770 1.150 ;
        RECT 333.310 0.770 333.690 1.150 ;
        RECT 333.970 0.770 334.350 1.150 ;
        RECT 334.630 0.770 335.010 1.150 ;
        RECT 335.550 0.770 335.930 1.150 ;
        RECT 336.210 0.770 336.590 1.150 ;
        RECT 336.870 0.770 337.250 1.150 ;
        RECT 337.790 0.770 338.170 1.150 ;
        RECT 338.450 0.770 338.830 1.150 ;
        RECT 339.110 0.770 339.490 1.150 ;
        RECT 340.030 0.770 340.410 1.150 ;
        RECT 340.690 0.770 341.070 1.150 ;
        RECT 341.350 0.770 341.730 1.150 ;
        RECT 342.390 0.770 342.770 1.150 ;
        RECT 343.390 0.770 343.770 1.150 ;
        RECT 344.050 0.770 344.430 1.150 ;
        RECT 344.710 0.770 345.090 1.150 ;
        RECT 345.630 0.770 346.010 1.150 ;
        RECT 346.290 0.770 346.670 1.150 ;
        RECT 346.950 0.770 347.330 1.150 ;
        RECT 347.870 0.770 348.250 1.150 ;
        RECT 348.530 0.770 348.910 1.150 ;
        RECT 349.190 0.770 349.570 1.150 ;
        RECT 350.110 0.770 350.490 1.150 ;
        RECT 350.770 0.770 351.150 1.150 ;
        RECT 351.430 0.770 351.810 1.150 ;
        RECT 352.190 0.770 352.570 1.150 ;
        RECT 353.510 0.770 353.890 1.150 ;
        RECT 355.710 0.770 356.090 1.150 ;
        RECT 356.370 0.770 356.750 1.150 ;
        RECT 357.030 0.770 357.410 1.150 ;
        RECT 357.950 0.770 358.330 1.150 ;
        RECT 358.610 0.770 358.990 1.150 ;
        RECT 359.270 0.770 359.650 1.150 ;
        RECT 360.190 0.770 360.570 1.150 ;
        RECT 360.850 0.770 361.230 1.150 ;
        RECT 361.510 0.770 361.890 1.150 ;
        RECT 362.550 0.770 362.930 1.150 ;
        RECT 363.550 0.770 363.930 1.150 ;
        RECT 364.210 0.770 364.590 1.150 ;
        RECT 364.870 0.770 365.250 1.150 ;
        RECT 365.790 0.770 366.170 1.150 ;
        RECT 366.450 0.770 366.830 1.150 ;
        RECT 367.110 0.770 367.490 1.150 ;
        RECT 368.030 0.770 368.410 1.150 ;
        RECT 368.690 0.770 369.070 1.150 ;
        RECT 369.350 0.770 369.730 1.150 ;
        RECT 370.270 0.770 370.650 1.150 ;
        RECT 370.930 0.770 371.310 1.150 ;
        RECT 371.590 0.770 371.970 1.150 ;
        RECT 372.510 0.770 372.890 1.150 ;
        RECT 373.170 0.770 373.550 1.150 ;
        RECT 373.830 0.770 374.210 1.150 ;
        RECT 374.750 0.770 375.130 1.150 ;
        RECT 375.410 0.770 375.790 1.150 ;
        RECT 376.070 0.770 376.450 1.150 ;
        RECT 376.990 0.770 377.370 1.150 ;
        RECT 377.650 0.770 378.030 1.150 ;
        RECT 378.310 0.770 378.690 1.150 ;
        RECT 379.230 0.770 379.610 1.150 ;
        RECT 379.890 0.770 380.270 1.150 ;
        RECT 380.550 0.770 380.930 1.150 ;
        RECT 381.470 0.770 381.850 1.150 ;
        RECT 382.130 0.770 382.510 1.150 ;
        RECT 382.790 0.770 383.170 1.150 ;
        RECT 383.830 0.770 384.210 1.150 ;
        RECT 384.830 0.770 385.210 1.150 ;
        RECT 385.490 0.770 385.870 1.150 ;
        RECT 386.150 0.770 386.530 1.150 ;
        RECT 387.070 0.770 387.450 1.150 ;
        RECT 387.730 0.770 388.110 1.150 ;
        RECT 388.390 0.770 388.770 1.150 ;
        RECT 389.310 0.770 389.690 1.150 ;
        RECT 389.970 0.770 390.350 1.150 ;
        RECT 390.630 0.770 391.010 1.150 ;
        RECT 391.550 0.770 391.930 1.150 ;
        RECT 392.210 0.770 392.590 1.150 ;
        RECT 392.870 0.770 393.250 1.150 ;
        RECT 393.790 0.770 394.170 1.150 ;
        RECT 394.450 0.770 394.830 1.150 ;
        RECT 395.110 0.770 395.490 1.150 ;
        RECT 395.870 0.770 396.250 1.150 ;
        RECT 397.190 0.770 397.570 1.150 ;
        RECT 399.390 0.770 399.770 1.150 ;
        RECT 400.050 0.770 400.430 1.150 ;
        RECT 400.710 0.770 401.090 1.150 ;
        RECT 401.630 0.770 402.010 1.150 ;
        RECT 402.290 0.770 402.670 1.150 ;
        RECT 402.950 0.770 403.330 1.150 ;
        RECT 403.990 0.770 404.370 1.150 ;
        RECT 404.990 0.770 405.370 1.150 ;
        RECT 405.650 0.770 406.030 1.150 ;
        RECT 406.310 0.770 406.690 1.150 ;
        RECT 407.230 0.770 407.610 1.150 ;
        RECT 407.890 0.770 408.270 1.150 ;
        RECT 408.550 0.770 408.930 1.150 ;
        RECT 409.470 0.770 409.850 1.150 ;
        RECT 410.130 0.770 410.510 1.150 ;
        RECT 410.790 0.770 411.170 1.150 ;
        RECT 411.710 0.770 412.090 1.150 ;
        RECT 412.370 0.770 412.750 1.150 ;
        RECT 413.030 0.770 413.410 1.150 ;
        RECT 413.950 0.770 414.330 1.150 ;
        RECT 414.610 0.770 414.990 1.150 ;
        RECT 415.270 0.770 415.650 1.150 ;
        RECT 416.190 0.770 416.570 1.150 ;
        RECT 416.850 0.770 417.230 1.150 ;
        RECT 417.510 0.770 417.890 1.150 ;
        RECT 418.430 0.770 418.810 1.150 ;
        RECT 419.090 0.770 419.470 1.150 ;
        RECT 419.750 0.770 420.130 1.150 ;
        RECT 420.670 0.770 421.050 1.150 ;
        RECT 421.330 0.770 421.710 1.150 ;
        RECT 421.990 0.770 422.370 1.150 ;
        RECT 422.910 0.770 423.290 1.150 ;
        RECT 423.570 0.770 423.950 1.150 ;
        RECT 424.230 0.770 424.610 1.150 ;
        RECT 425.270 0.770 425.650 1.150 ;
        RECT 426.270 0.770 426.650 1.150 ;
        RECT 426.930 0.770 427.310 1.150 ;
        RECT 427.590 0.770 427.970 1.150 ;
        RECT 428.510 0.770 428.890 1.150 ;
        RECT 429.170 0.770 429.550 1.150 ;
        RECT 429.830 0.770 430.210 1.150 ;
        RECT 430.750 0.770 431.130 1.150 ;
        RECT 431.410 0.770 431.790 1.150 ;
        RECT 432.070 0.770 432.450 1.150 ;
        RECT 432.990 0.770 433.370 1.150 ;
        RECT 433.650 0.770 434.030 1.150 ;
        RECT 434.310 0.770 434.690 1.150 ;
        RECT 435.230 0.770 435.610 1.150 ;
        RECT 435.890 0.770 436.270 1.150 ;
        RECT 436.550 0.770 436.930 1.150 ;
        RECT 437.310 0.770 437.690 1.150 ;
        RECT 438.630 0.770 439.010 1.150 ;
        RECT 440.830 0.770 441.210 1.150 ;
        RECT 441.490 0.770 441.870 1.150 ;
        RECT 442.150 0.770 442.530 1.150 ;
        RECT 443.070 0.770 443.450 1.150 ;
        RECT 443.730 0.770 444.110 1.150 ;
        RECT 444.390 0.770 444.770 1.150 ;
        RECT 445.430 0.770 445.810 1.150 ;
        RECT 446.430 0.770 446.810 1.150 ;
        RECT 447.090 0.770 447.470 1.150 ;
        RECT 447.750 0.770 448.130 1.150 ;
        RECT 448.670 0.770 449.050 1.150 ;
        RECT 449.330 0.770 449.710 1.150 ;
        RECT 449.990 0.770 450.370 1.150 ;
        RECT 450.910 0.770 451.290 1.150 ;
        RECT 451.570 0.770 451.950 1.150 ;
        RECT 452.230 0.770 452.610 1.150 ;
        RECT 453.150 0.770 453.530 1.150 ;
        RECT 453.810 0.770 454.190 1.150 ;
        RECT 454.470 0.770 454.850 1.150 ;
        RECT 455.390 0.770 455.770 1.150 ;
        RECT 456.050 0.770 456.430 1.150 ;
        RECT 456.710 0.770 457.090 1.150 ;
        RECT 457.630 0.770 458.010 1.150 ;
        RECT 458.290 0.770 458.670 1.150 ;
        RECT 458.950 0.770 459.330 1.150 ;
        RECT 459.870 0.770 460.250 1.150 ;
        RECT 460.530 0.770 460.910 1.150 ;
        RECT 461.190 0.770 461.570 1.150 ;
        RECT 462.110 0.770 462.490 1.150 ;
        RECT 462.770 0.770 463.150 1.150 ;
        RECT 463.430 0.770 463.810 1.150 ;
        RECT 464.350 0.770 464.730 1.150 ;
        RECT 465.010 0.770 465.390 1.150 ;
        RECT 465.670 0.770 466.050 1.150 ;
        RECT 466.710 0.770 467.090 1.150 ;
        RECT 467.710 0.770 468.090 1.150 ;
        RECT 468.370 0.770 468.750 1.150 ;
        RECT 469.030 0.770 469.410 1.150 ;
        RECT 469.950 0.770 470.330 1.150 ;
        RECT 470.610 0.770 470.990 1.150 ;
        RECT 471.270 0.770 471.650 1.150 ;
        RECT 472.190 0.770 472.570 1.150 ;
        RECT 472.850 0.770 473.230 1.150 ;
        RECT 473.510 0.770 473.890 1.150 ;
        RECT 474.430 0.770 474.810 1.150 ;
        RECT 475.090 0.770 475.470 1.150 ;
        RECT 475.750 0.770 476.130 1.150 ;
        RECT 476.670 0.770 477.050 1.150 ;
        RECT 477.330 0.770 477.710 1.150 ;
        RECT 477.990 0.770 478.370 1.150 ;
        RECT 478.910 0.770 479.290 1.150 ;
        RECT 479.570 0.770 479.950 1.150 ;
        RECT 480.230 0.770 480.610 1.150 ;
        RECT 480.990 0.770 481.370 1.150 ;
        RECT 482.310 0.770 482.690 1.150 ;
        RECT 484.510 0.770 484.890 1.150 ;
        RECT 485.170 0.770 485.550 1.150 ;
        RECT 485.830 0.770 486.210 1.150 ;
        RECT 486.870 0.770 487.250 1.150 ;
        RECT 487.870 0.770 488.250 1.150 ;
        RECT 488.530 0.770 488.910 1.150 ;
        RECT 489.190 0.770 489.570 1.150 ;
        RECT 490.110 0.770 490.490 1.150 ;
        RECT 490.770 0.770 491.150 1.150 ;
        RECT 491.430 0.770 491.810 1.150 ;
        RECT 492.350 0.770 492.730 1.150 ;
        RECT 493.010 0.770 493.390 1.150 ;
        RECT 493.670 0.770 494.050 1.150 ;
        RECT 494.590 0.770 494.970 1.150 ;
        RECT 495.250 0.770 495.630 1.150 ;
        RECT 495.910 0.770 496.290 1.150 ;
        RECT 496.830 0.770 497.210 1.150 ;
        RECT 497.490 0.770 497.870 1.150 ;
        RECT 498.150 0.770 498.530 1.150 ;
        RECT 499.070 0.770 499.450 1.150 ;
        RECT 499.730 0.770 500.110 1.150 ;
        RECT 500.390 0.770 500.770 1.150 ;
        RECT 501.310 0.770 501.690 1.150 ;
        RECT 501.970 0.770 502.350 1.150 ;
        RECT 502.630 0.770 503.010 1.150 ;
        RECT 503.550 0.770 503.930 1.150 ;
        RECT 504.210 0.770 504.590 1.150 ;
        RECT 504.870 0.770 505.250 1.150 ;
        RECT 505.790 0.770 506.170 1.150 ;
        RECT 506.450 0.770 506.830 1.150 ;
        RECT 507.110 0.770 507.490 1.150 ;
        RECT 508.150 0.770 508.530 1.150 ;
        RECT 509.150 0.770 509.530 1.150 ;
        RECT 509.810 0.770 510.190 1.150 ;
        RECT 510.470 0.770 510.850 1.150 ;
        RECT 511.390 0.770 511.770 1.150 ;
        RECT 512.050 0.770 512.430 1.150 ;
        RECT 512.710 0.770 513.090 1.150 ;
        RECT 513.630 0.770 514.010 1.150 ;
        RECT 514.290 0.770 514.670 1.150 ;
        RECT 514.950 0.770 515.330 1.150 ;
        RECT 515.870 0.770 516.250 1.150 ;
        RECT 516.530 0.770 516.910 1.150 ;
        RECT 517.190 0.770 517.570 1.150 ;
        RECT 518.110 0.770 518.490 1.150 ;
        RECT 518.770 0.770 519.150 1.150 ;
        RECT 519.430 0.770 519.810 1.150 ;
        RECT 520.350 0.770 520.730 1.150 ;
        RECT 521.010 0.770 521.390 1.150 ;
        RECT 521.670 0.770 522.050 1.150 ;
        RECT 522.430 0.770 522.810 1.150 ;
        RECT 523.750 0.770 524.130 1.150 ;
        RECT 525.950 0.770 526.330 1.150 ;
        RECT 526.610 0.770 526.990 1.150 ;
        RECT 527.270 0.770 527.650 1.150 ;
        RECT 528.310 0.770 528.690 1.150 ;
        RECT 529.310 0.770 529.690 1.150 ;
        RECT 529.970 0.770 530.350 1.150 ;
        RECT 530.630 0.770 531.010 1.150 ;
        RECT 531.550 0.770 531.930 1.150 ;
        RECT 532.210 0.770 532.590 1.150 ;
        RECT 532.870 0.770 533.250 1.150 ;
        RECT 533.790 0.770 534.170 1.150 ;
        RECT 534.450 0.770 534.830 1.150 ;
        RECT 535.110 0.770 535.490 1.150 ;
        RECT 536.030 0.770 536.410 1.150 ;
        RECT 536.690 0.770 537.070 1.150 ;
        RECT 537.350 0.770 537.730 1.150 ;
        RECT 538.270 0.770 538.650 1.150 ;
        RECT 538.930 0.770 539.310 1.150 ;
        RECT 539.590 0.770 539.970 1.150 ;
        RECT 540.510 0.770 540.890 1.150 ;
        RECT 541.170 0.770 541.550 1.150 ;
        RECT 541.830 0.770 542.210 1.150 ;
        RECT 542.750 0.770 543.130 1.150 ;
        RECT 543.410 0.770 543.790 1.150 ;
        RECT 544.070 0.770 544.450 1.150 ;
        RECT 544.990 0.770 545.370 1.150 ;
        RECT 545.650 0.770 546.030 1.150 ;
        RECT 546.310 0.770 546.690 1.150 ;
        RECT 547.230 0.770 547.610 1.150 ;
        RECT 547.890 0.770 548.270 1.150 ;
        RECT 548.550 0.770 548.930 1.150 ;
        RECT 549.590 0.770 549.970 1.150 ;
        RECT 550.590 0.770 550.970 1.150 ;
        RECT 551.250 0.770 551.630 1.150 ;
        RECT 551.910 0.770 552.290 1.150 ;
        RECT 552.830 0.770 553.210 1.150 ;
        RECT 553.490 0.770 553.870 1.150 ;
        RECT 554.150 0.770 554.530 1.150 ;
        RECT 555.070 0.770 555.450 1.150 ;
        RECT 555.730 0.770 556.110 1.150 ;
        RECT 556.390 0.770 556.770 1.150 ;
        RECT 557.310 0.770 557.690 1.150 ;
        RECT 557.970 0.770 558.350 1.150 ;
        RECT 558.630 0.770 559.010 1.150 ;
        RECT 559.550 0.770 559.930 1.150 ;
        RECT 560.210 0.770 560.590 1.150 ;
        RECT 560.870 0.770 561.250 1.150 ;
        RECT 561.790 0.770 562.170 1.150 ;
        RECT 562.450 0.770 562.830 1.150 ;
        RECT 563.110 0.770 563.490 1.150 ;
        RECT 564.030 0.770 564.410 1.150 ;
        RECT 564.690 0.770 565.070 1.150 ;
        RECT 565.350 0.770 565.730 1.150 ;
        RECT 566.110 0.770 566.490 1.150 ;
        RECT 567.430 0.770 567.810 1.150 ;
        RECT 569.750 0.770 570.130 1.150 ;
        RECT 570.750 0.770 571.130 1.150 ;
        RECT 571.410 0.770 571.790 1.150 ;
        RECT 572.070 0.770 572.450 1.150 ;
        RECT 572.990 0.770 573.370 1.150 ;
        RECT 573.650 0.770 574.030 1.150 ;
        RECT 574.310 0.770 574.690 1.150 ;
        RECT 575.230 0.770 575.610 1.150 ;
        RECT 575.890 0.770 576.270 1.150 ;
        RECT 576.550 0.770 576.930 1.150 ;
        RECT 577.470 0.770 577.850 1.150 ;
        RECT 578.130 0.770 578.510 1.150 ;
        RECT 578.790 0.770 579.170 1.150 ;
        RECT 579.710 0.770 580.090 1.150 ;
        RECT 580.370 0.770 580.750 1.150 ;
        RECT 581.030 0.770 581.410 1.150 ;
        RECT 581.950 0.770 582.330 1.150 ;
        RECT 582.610 0.770 582.990 1.150 ;
        RECT 583.270 0.770 583.650 1.150 ;
        RECT 584.190 0.770 584.570 1.150 ;
        RECT 584.850 0.770 585.230 1.150 ;
        RECT 585.510 0.770 585.890 1.150 ;
        RECT 586.430 0.770 586.810 1.150 ;
        RECT 587.090 0.770 587.470 1.150 ;
        RECT 587.750 0.770 588.130 1.150 ;
        RECT 588.670 0.770 589.050 1.150 ;
        RECT 589.330 0.770 589.710 1.150 ;
        RECT 589.990 0.770 590.370 1.150 ;
        RECT 591.030 0.770 591.410 1.150 ;
        RECT 592.030 0.770 592.410 1.150 ;
        RECT 592.690 0.770 593.070 1.150 ;
        RECT 593.350 0.770 593.730 1.150 ;
        RECT 594.270 0.770 594.650 1.150 ;
        RECT 594.930 0.770 595.310 1.150 ;
        RECT 595.590 0.770 595.970 1.150 ;
        RECT 596.510 0.770 596.890 1.150 ;
        RECT 597.170 0.770 597.550 1.150 ;
        RECT 597.830 0.770 598.210 1.150 ;
        RECT 598.750 0.770 599.130 1.150 ;
        RECT 599.410 0.770 599.790 1.150 ;
        RECT 600.070 0.770 600.450 1.150 ;
        RECT 600.990 0.770 601.370 1.150 ;
        RECT 601.650 0.770 602.030 1.150 ;
        RECT 602.310 0.770 602.690 1.150 ;
        RECT 603.230 0.770 603.610 1.150 ;
        RECT 603.890 0.770 604.270 1.150 ;
        RECT 604.550 0.770 604.930 1.150 ;
        RECT 605.470 0.770 605.850 1.150 ;
        RECT 606.130 0.770 606.510 1.150 ;
        RECT 606.790 0.770 607.170 1.150 ;
        RECT 607.550 0.770 607.930 1.150 ;
        RECT 608.870 0.770 609.250 1.150 ;
        RECT 611.190 0.770 611.570 1.150 ;
        RECT 612.190 0.770 612.570 1.150 ;
        RECT 612.850 0.770 613.230 1.150 ;
        RECT 613.510 0.770 613.890 1.150 ;
        RECT 614.430 0.770 614.810 1.150 ;
        RECT 615.090 0.770 615.470 1.150 ;
        RECT 615.750 0.770 616.130 1.150 ;
        RECT 616.670 0.770 617.050 1.150 ;
        RECT 617.330 0.770 617.710 1.150 ;
        RECT 617.990 0.770 618.370 1.150 ;
        RECT 618.910 0.770 619.290 1.150 ;
        RECT 619.570 0.770 619.950 1.150 ;
        RECT 620.230 0.770 620.610 1.150 ;
        RECT 621.150 0.770 621.530 1.150 ;
        RECT 621.810 0.770 622.190 1.150 ;
        RECT 622.470 0.770 622.850 1.150 ;
        RECT 623.390 0.770 623.770 1.150 ;
        RECT 624.050 0.770 624.430 1.150 ;
        RECT 624.710 0.770 625.090 1.150 ;
        RECT 625.630 0.770 626.010 1.150 ;
        RECT 626.290 0.770 626.670 1.150 ;
        RECT 626.950 0.770 627.330 1.150 ;
        RECT 627.870 0.770 628.250 1.150 ;
        RECT 628.530 0.770 628.910 1.150 ;
        RECT 629.190 0.770 629.570 1.150 ;
        RECT 630.110 0.770 630.490 1.150 ;
        RECT 630.770 0.770 631.150 1.150 ;
        RECT 631.430 0.770 631.810 1.150 ;
        RECT 632.470 0.770 632.850 1.150 ;
        RECT 633.470 0.770 633.850 1.150 ;
        RECT 634.130 0.770 634.510 1.150 ;
        RECT 634.790 0.770 635.170 1.150 ;
        RECT 635.710 0.770 636.090 1.150 ;
        RECT 636.370 0.770 636.750 1.150 ;
        RECT 637.030 0.770 637.410 1.150 ;
        RECT 637.950 0.770 638.330 1.150 ;
        RECT 638.610 0.770 638.990 1.150 ;
        RECT 639.270 0.770 639.650 1.150 ;
        RECT 640.190 0.770 640.570 1.150 ;
        RECT 640.850 0.770 641.230 1.150 ;
        RECT 641.510 0.770 641.890 1.150 ;
        RECT 642.430 0.770 642.810 1.150 ;
        RECT 643.090 0.770 643.470 1.150 ;
        RECT 643.750 0.770 644.130 1.150 ;
        RECT 644.670 0.770 645.050 1.150 ;
        RECT 645.330 0.770 645.710 1.150 ;
        RECT 645.990 0.770 646.370 1.150 ;
        RECT 646.910 0.770 647.290 1.150 ;
        RECT 647.570 0.770 647.950 1.150 ;
        RECT 648.230 0.770 648.610 1.150 ;
        RECT 649.150 0.770 649.530 1.150 ;
        RECT 649.810 0.770 650.190 1.150 ;
        RECT 650.470 0.770 650.850 1.150 ;
        RECT 651.230 0.770 651.610 1.150 ;
        RECT 652.550 0.770 652.930 1.150 ;
        RECT 654.870 0.770 655.250 1.150 ;
        RECT 655.870 0.770 656.250 1.150 ;
        RECT 656.530 0.770 656.910 1.150 ;
        RECT 657.190 0.770 657.570 1.150 ;
        RECT 658.110 0.770 658.490 1.150 ;
        RECT 658.770 0.770 659.150 1.150 ;
        RECT 659.430 0.770 659.810 1.150 ;
        RECT 660.350 0.770 660.730 1.150 ;
        RECT 661.010 0.770 661.390 1.150 ;
        RECT 661.670 0.770 662.050 1.150 ;
        RECT 662.590 0.770 662.970 1.150 ;
        RECT 663.250 0.770 663.630 1.150 ;
        RECT 663.910 0.770 664.290 1.150 ;
        RECT 664.830 0.770 665.210 1.150 ;
        RECT 665.490 0.770 665.870 1.150 ;
        RECT 666.150 0.770 666.530 1.150 ;
        RECT 667.070 0.770 667.450 1.150 ;
        RECT 667.730 0.770 668.110 1.150 ;
        RECT 668.390 0.770 668.770 1.150 ;
        RECT 669.310 0.770 669.690 1.150 ;
        RECT 669.970 0.770 670.350 1.150 ;
        RECT 670.630 0.770 671.010 1.150 ;
        RECT 671.550 0.770 671.930 1.150 ;
        RECT 672.210 0.770 672.590 1.150 ;
        RECT 672.870 0.770 673.250 1.150 ;
        RECT 673.790 0.770 674.170 1.150 ;
        RECT 674.450 0.770 674.830 1.150 ;
        RECT 675.110 0.770 675.490 1.150 ;
        RECT 676.150 0.770 676.530 1.150 ;
        RECT 677.150 0.770 677.530 1.150 ;
        RECT 677.810 0.770 678.190 1.150 ;
        RECT 678.470 0.770 678.850 1.150 ;
        RECT 679.490 0.770 679.870 1.150 ;
      LAYER Via2 ;
        RECT 0.815 58.795 1.095 59.075 ;
        RECT 0.815 58.135 1.095 58.415 ;
        RECT 0.815 57.475 1.095 57.755 ;
        RECT 0.815 56.815 1.095 57.095 ;
        RECT 0.815 56.155 1.095 56.435 ;
        RECT 0.815 55.495 1.095 55.775 ;
        RECT 0.815 54.835 1.095 55.115 ;
        RECT 0.815 54.175 1.095 54.455 ;
        RECT 0.815 53.515 1.095 53.795 ;
        RECT 0.815 52.855 1.095 53.135 ;
        RECT 0.815 52.195 1.095 52.475 ;
        RECT 0.815 51.535 1.095 51.815 ;
        RECT 0.815 50.875 1.095 51.155 ;
        RECT 0.815 50.215 1.095 50.495 ;
        RECT 5.300 47.855 5.580 48.135 ;
        RECT 5.960 47.855 6.240 48.135 ;
        RECT 6.620 47.855 6.900 48.135 ;
        RECT 5.300 47.195 5.580 47.475 ;
        RECT 5.960 47.195 6.240 47.475 ;
        RECT 6.620 47.195 6.900 47.475 ;
        RECT 5.300 46.535 5.580 46.815 ;
        RECT 5.960 46.535 6.240 46.815 ;
        RECT 6.620 46.535 6.900 46.815 ;
        RECT 5.300 22.255 5.580 22.535 ;
        RECT 5.960 22.255 6.240 22.535 ;
        RECT 6.620 22.255 6.900 22.535 ;
        RECT 5.300 21.595 5.580 21.875 ;
        RECT 5.960 21.595 6.240 21.875 ;
        RECT 6.620 21.595 6.900 21.875 ;
        RECT 5.300 20.935 5.580 21.215 ;
        RECT 5.960 20.935 6.240 21.215 ;
        RECT 6.620 20.935 6.900 21.215 ;
        RECT 11.105 58.795 11.385 59.075 ;
        RECT 11.105 58.135 11.385 58.415 ;
        RECT 11.105 57.475 11.385 57.755 ;
        RECT 11.105 56.815 11.385 57.095 ;
        RECT 11.105 56.155 11.385 56.435 ;
        RECT 11.105 55.495 11.385 55.775 ;
        RECT 11.105 54.835 11.385 55.115 ;
        RECT 11.105 54.175 11.385 54.455 ;
        RECT 11.105 53.515 11.385 53.795 ;
        RECT 11.105 52.855 11.385 53.135 ;
        RECT 11.105 52.195 11.385 52.475 ;
        RECT 11.105 51.535 11.385 51.815 ;
        RECT 11.105 50.875 11.385 51.155 ;
        RECT 11.105 50.215 11.385 50.495 ;
        RECT 21.390 58.795 21.670 59.075 ;
        RECT 21.390 58.135 21.670 58.415 ;
        RECT 21.390 57.475 21.670 57.755 ;
        RECT 21.390 56.815 21.670 57.095 ;
        RECT 21.390 56.155 21.670 56.435 ;
        RECT 21.390 55.495 21.670 55.775 ;
        RECT 21.390 54.835 21.670 55.115 ;
        RECT 21.390 54.175 21.670 54.455 ;
        RECT 21.390 53.515 21.670 53.795 ;
        RECT 21.390 52.855 21.670 53.135 ;
        RECT 21.390 52.195 21.670 52.475 ;
        RECT 21.390 51.535 21.670 51.815 ;
        RECT 21.390 50.875 21.670 51.155 ;
        RECT 21.390 50.215 21.670 50.495 ;
        RECT 15.600 45.155 15.880 45.435 ;
        RECT 16.260 45.155 16.540 45.435 ;
        RECT 16.920 45.155 17.200 45.435 ;
        RECT 15.600 44.495 15.880 44.775 ;
        RECT 16.260 44.495 16.540 44.775 ;
        RECT 16.920 44.495 17.200 44.775 ;
        RECT 15.600 43.835 15.880 44.115 ;
        RECT 16.260 43.835 16.540 44.115 ;
        RECT 16.920 43.835 17.200 44.115 ;
        RECT 25.875 42.455 26.155 42.735 ;
        RECT 26.535 42.455 26.815 42.735 ;
        RECT 27.195 42.455 27.475 42.735 ;
        RECT 25.875 41.795 26.155 42.075 ;
        RECT 26.535 41.795 26.815 42.075 ;
        RECT 27.195 41.795 27.475 42.075 ;
        RECT 25.875 41.135 26.155 41.415 ;
        RECT 26.535 41.135 26.815 41.415 ;
        RECT 27.195 41.135 27.475 41.415 ;
        RECT 25.875 27.655 26.155 27.935 ;
        RECT 26.535 27.655 26.815 27.935 ;
        RECT 27.195 27.655 27.475 27.935 ;
        RECT 25.875 26.995 26.155 27.275 ;
        RECT 26.535 26.995 26.815 27.275 ;
        RECT 27.195 26.995 27.475 27.275 ;
        RECT 25.875 26.335 26.155 26.615 ;
        RECT 26.535 26.335 26.815 26.615 ;
        RECT 27.195 26.335 27.475 26.615 ;
        RECT 15.600 24.955 15.880 25.235 ;
        RECT 16.260 24.955 16.540 25.235 ;
        RECT 16.920 24.955 17.200 25.235 ;
        RECT 15.600 24.295 15.880 24.575 ;
        RECT 16.260 24.295 16.540 24.575 ;
        RECT 16.920 24.295 17.200 24.575 ;
        RECT 15.600 23.635 15.880 23.915 ;
        RECT 16.260 23.635 16.540 23.915 ;
        RECT 16.920 23.635 17.200 23.915 ;
        RECT 31.680 58.795 31.960 59.075 ;
        RECT 31.680 58.135 31.960 58.415 ;
        RECT 31.680 57.475 31.960 57.755 ;
        RECT 31.680 56.815 31.960 57.095 ;
        RECT 31.680 56.155 31.960 56.435 ;
        RECT 31.680 55.495 31.960 55.775 ;
        RECT 31.680 54.835 31.960 55.115 ;
        RECT 31.680 54.175 31.960 54.455 ;
        RECT 31.680 53.515 31.960 53.795 ;
        RECT 31.680 52.855 31.960 53.135 ;
        RECT 31.680 52.195 31.960 52.475 ;
        RECT 31.680 51.535 31.960 51.815 ;
        RECT 31.680 50.875 31.960 51.155 ;
        RECT 31.680 50.215 31.960 50.495 ;
        RECT 41.965 58.795 42.245 59.075 ;
        RECT 43.385 58.795 43.665 59.075 ;
        RECT 41.965 58.135 42.245 58.415 ;
        RECT 43.385 58.135 43.665 58.415 ;
        RECT 41.965 57.475 42.245 57.755 ;
        RECT 43.385 57.475 43.665 57.755 ;
        RECT 41.965 56.815 42.245 57.095 ;
        RECT 43.385 56.815 43.665 57.095 ;
        RECT 41.965 56.155 42.245 56.435 ;
        RECT 43.385 56.155 43.665 56.435 ;
        RECT 41.965 55.495 42.245 55.775 ;
        RECT 43.385 55.495 43.665 55.775 ;
        RECT 41.965 54.835 42.245 55.115 ;
        RECT 43.385 54.835 43.665 55.115 ;
        RECT 41.965 54.175 42.245 54.455 ;
        RECT 43.385 54.175 43.665 54.455 ;
        RECT 41.965 53.515 42.245 53.795 ;
        RECT 43.385 53.515 43.665 53.795 ;
        RECT 41.965 52.855 42.245 53.135 ;
        RECT 43.385 52.855 43.665 53.135 ;
        RECT 41.965 52.195 42.245 52.475 ;
        RECT 43.385 52.195 43.665 52.475 ;
        RECT 41.965 51.535 42.245 51.815 ;
        RECT 43.385 51.535 43.665 51.815 ;
        RECT 41.965 50.875 42.245 51.155 ;
        RECT 43.385 50.875 43.665 51.155 ;
        RECT 41.965 50.215 42.245 50.495 ;
        RECT 43.385 50.215 43.665 50.495 ;
        RECT 47.870 47.855 48.150 48.135 ;
        RECT 48.530 47.855 48.810 48.135 ;
        RECT 49.190 47.855 49.470 48.135 ;
        RECT 47.870 47.195 48.150 47.475 ;
        RECT 48.530 47.195 48.810 47.475 ;
        RECT 49.190 47.195 49.470 47.475 ;
        RECT 47.870 46.535 48.150 46.815 ;
        RECT 48.530 46.535 48.810 46.815 ;
        RECT 49.190 46.535 49.470 46.815 ;
        RECT 36.175 39.755 36.455 40.035 ;
        RECT 36.835 39.755 37.115 40.035 ;
        RECT 37.495 39.755 37.775 40.035 ;
        RECT 36.175 39.095 36.455 39.375 ;
        RECT 36.835 39.095 37.115 39.375 ;
        RECT 37.495 39.095 37.775 39.375 ;
        RECT 36.175 38.435 36.455 38.715 ;
        RECT 36.835 38.435 37.115 38.715 ;
        RECT 37.495 38.435 37.775 38.715 ;
        RECT 36.175 30.355 36.455 30.635 ;
        RECT 36.835 30.355 37.115 30.635 ;
        RECT 37.495 30.355 37.775 30.635 ;
        RECT 36.175 29.695 36.455 29.975 ;
        RECT 36.835 29.695 37.115 29.975 ;
        RECT 37.495 29.695 37.775 29.975 ;
        RECT 36.175 29.035 36.455 29.315 ;
        RECT 36.835 29.035 37.115 29.315 ;
        RECT 37.495 29.035 37.775 29.315 ;
        RECT 47.870 22.255 48.150 22.535 ;
        RECT 48.530 22.255 48.810 22.535 ;
        RECT 49.190 22.255 49.470 22.535 ;
        RECT 47.870 21.595 48.150 21.875 ;
        RECT 48.530 21.595 48.810 21.875 ;
        RECT 49.190 21.595 49.470 21.875 ;
        RECT 47.870 20.935 48.150 21.215 ;
        RECT 48.530 20.935 48.810 21.215 ;
        RECT 49.190 20.935 49.470 21.215 ;
        RECT 4.660 8.140 4.940 8.420 ;
        RECT 4.660 7.480 4.940 7.760 ;
        RECT 4.660 6.820 4.940 7.100 ;
        RECT 0.900 4.740 1.180 5.020 ;
        RECT 2.040 4.740 2.320 5.020 ;
        RECT 8.080 4.770 8.360 5.050 ;
        RECT 8.740 4.770 9.020 5.050 ;
        RECT 9.400 4.770 9.680 5.050 ;
        RECT 14.610 4.740 14.890 5.020 ;
        RECT 15.270 4.740 15.550 5.020 ;
        RECT 15.930 4.740 16.210 5.020 ;
        RECT 17.970 4.740 18.250 5.020 ;
        RECT 18.630 4.740 18.910 5.020 ;
        RECT 19.290 4.740 19.570 5.020 ;
        RECT 53.675 58.795 53.955 59.075 ;
        RECT 53.675 58.135 53.955 58.415 ;
        RECT 53.675 57.475 53.955 57.755 ;
        RECT 53.675 56.815 53.955 57.095 ;
        RECT 53.675 56.155 53.955 56.435 ;
        RECT 53.675 55.495 53.955 55.775 ;
        RECT 53.675 54.835 53.955 55.115 ;
        RECT 53.675 54.175 53.955 54.455 ;
        RECT 53.675 53.515 53.955 53.795 ;
        RECT 53.675 52.855 53.955 53.135 ;
        RECT 53.675 52.195 53.955 52.475 ;
        RECT 53.675 51.535 53.955 51.815 ;
        RECT 53.675 50.875 53.955 51.155 ;
        RECT 53.675 50.215 53.955 50.495 ;
        RECT 63.960 58.795 64.240 59.075 ;
        RECT 63.960 58.135 64.240 58.415 ;
        RECT 63.960 57.475 64.240 57.755 ;
        RECT 63.960 56.815 64.240 57.095 ;
        RECT 63.960 56.155 64.240 56.435 ;
        RECT 63.960 55.495 64.240 55.775 ;
        RECT 63.960 54.835 64.240 55.115 ;
        RECT 63.960 54.175 64.240 54.455 ;
        RECT 63.960 53.515 64.240 53.795 ;
        RECT 63.960 52.855 64.240 53.135 ;
        RECT 63.960 52.195 64.240 52.475 ;
        RECT 63.960 51.535 64.240 51.815 ;
        RECT 63.960 50.875 64.240 51.155 ;
        RECT 63.960 50.215 64.240 50.495 ;
        RECT 58.170 45.155 58.450 45.435 ;
        RECT 58.830 45.155 59.110 45.435 ;
        RECT 59.490 45.155 59.770 45.435 ;
        RECT 58.170 44.495 58.450 44.775 ;
        RECT 58.830 44.495 59.110 44.775 ;
        RECT 59.490 44.495 59.770 44.775 ;
        RECT 58.170 43.835 58.450 44.115 ;
        RECT 58.830 43.835 59.110 44.115 ;
        RECT 59.490 43.835 59.770 44.115 ;
        RECT 68.445 42.455 68.725 42.735 ;
        RECT 69.105 42.455 69.385 42.735 ;
        RECT 69.765 42.455 70.045 42.735 ;
        RECT 68.445 41.795 68.725 42.075 ;
        RECT 69.105 41.795 69.385 42.075 ;
        RECT 69.765 41.795 70.045 42.075 ;
        RECT 68.445 41.135 68.725 41.415 ;
        RECT 69.105 41.135 69.385 41.415 ;
        RECT 69.765 41.135 70.045 41.415 ;
        RECT 68.445 27.655 68.725 27.935 ;
        RECT 69.105 27.655 69.385 27.935 ;
        RECT 69.765 27.655 70.045 27.935 ;
        RECT 68.445 26.995 68.725 27.275 ;
        RECT 69.105 26.995 69.385 27.275 ;
        RECT 69.765 26.995 70.045 27.275 ;
        RECT 68.445 26.335 68.725 26.615 ;
        RECT 69.105 26.335 69.385 26.615 ;
        RECT 69.765 26.335 70.045 26.615 ;
        RECT 58.170 24.955 58.450 25.235 ;
        RECT 58.830 24.955 59.110 25.235 ;
        RECT 59.490 24.955 59.770 25.235 ;
        RECT 58.170 24.295 58.450 24.575 ;
        RECT 58.830 24.295 59.110 24.575 ;
        RECT 59.490 24.295 59.770 24.575 ;
        RECT 58.170 23.635 58.450 23.915 ;
        RECT 58.830 23.635 59.110 23.915 ;
        RECT 59.490 23.635 59.770 23.915 ;
        RECT 74.250 58.795 74.530 59.075 ;
        RECT 74.250 58.135 74.530 58.415 ;
        RECT 74.250 57.475 74.530 57.755 ;
        RECT 74.250 56.815 74.530 57.095 ;
        RECT 74.250 56.155 74.530 56.435 ;
        RECT 74.250 55.495 74.530 55.775 ;
        RECT 74.250 54.835 74.530 55.115 ;
        RECT 74.250 54.175 74.530 54.455 ;
        RECT 74.250 53.515 74.530 53.795 ;
        RECT 74.250 52.855 74.530 53.135 ;
        RECT 74.250 52.195 74.530 52.475 ;
        RECT 74.250 51.535 74.530 51.815 ;
        RECT 74.250 50.875 74.530 51.155 ;
        RECT 74.250 50.215 74.530 50.495 ;
        RECT 84.535 58.795 84.815 59.075 ;
        RECT 85.955 58.795 86.235 59.075 ;
        RECT 84.535 58.135 84.815 58.415 ;
        RECT 85.955 58.135 86.235 58.415 ;
        RECT 84.535 57.475 84.815 57.755 ;
        RECT 85.955 57.475 86.235 57.755 ;
        RECT 84.535 56.815 84.815 57.095 ;
        RECT 85.955 56.815 86.235 57.095 ;
        RECT 84.535 56.155 84.815 56.435 ;
        RECT 85.955 56.155 86.235 56.435 ;
        RECT 84.535 55.495 84.815 55.775 ;
        RECT 85.955 55.495 86.235 55.775 ;
        RECT 84.535 54.835 84.815 55.115 ;
        RECT 85.955 54.835 86.235 55.115 ;
        RECT 84.535 54.175 84.815 54.455 ;
        RECT 85.955 54.175 86.235 54.455 ;
        RECT 84.535 53.515 84.815 53.795 ;
        RECT 85.955 53.515 86.235 53.795 ;
        RECT 84.535 52.855 84.815 53.135 ;
        RECT 85.955 52.855 86.235 53.135 ;
        RECT 84.535 52.195 84.815 52.475 ;
        RECT 85.955 52.195 86.235 52.475 ;
        RECT 84.535 51.535 84.815 51.815 ;
        RECT 85.955 51.535 86.235 51.815 ;
        RECT 84.535 50.875 84.815 51.155 ;
        RECT 85.955 50.875 86.235 51.155 ;
        RECT 84.535 50.215 84.815 50.495 ;
        RECT 85.955 50.215 86.235 50.495 ;
        RECT 90.440 47.855 90.720 48.135 ;
        RECT 91.100 47.855 91.380 48.135 ;
        RECT 91.760 47.855 92.040 48.135 ;
        RECT 90.440 47.195 90.720 47.475 ;
        RECT 91.100 47.195 91.380 47.475 ;
        RECT 91.760 47.195 92.040 47.475 ;
        RECT 90.440 46.535 90.720 46.815 ;
        RECT 91.100 46.535 91.380 46.815 ;
        RECT 91.760 46.535 92.040 46.815 ;
        RECT 78.745 39.755 79.025 40.035 ;
        RECT 79.405 39.755 79.685 40.035 ;
        RECT 80.065 39.755 80.345 40.035 ;
        RECT 78.745 39.095 79.025 39.375 ;
        RECT 79.405 39.095 79.685 39.375 ;
        RECT 80.065 39.095 80.345 39.375 ;
        RECT 78.745 38.435 79.025 38.715 ;
        RECT 79.405 38.435 79.685 38.715 ;
        RECT 80.065 38.435 80.345 38.715 ;
        RECT 78.745 30.355 79.025 30.635 ;
        RECT 79.405 30.355 79.685 30.635 ;
        RECT 80.065 30.355 80.345 30.635 ;
        RECT 78.745 29.695 79.025 29.975 ;
        RECT 79.405 29.695 79.685 29.975 ;
        RECT 80.065 29.695 80.345 29.975 ;
        RECT 78.745 29.035 79.025 29.315 ;
        RECT 79.405 29.035 79.685 29.315 ;
        RECT 80.065 29.035 80.345 29.315 ;
        RECT 90.440 22.255 90.720 22.535 ;
        RECT 91.100 22.255 91.380 22.535 ;
        RECT 91.760 22.255 92.040 22.535 ;
        RECT 90.440 21.595 90.720 21.875 ;
        RECT 91.100 21.595 91.380 21.875 ;
        RECT 91.760 21.595 92.040 21.875 ;
        RECT 90.440 20.935 90.720 21.215 ;
        RECT 91.100 20.935 91.380 21.215 ;
        RECT 91.760 20.935 92.040 21.215 ;
        RECT 22.850 8.140 23.130 8.420 ;
        RECT 38.800 8.140 39.080 8.420 ;
        RECT 53.630 8.140 53.910 8.420 ;
        RECT 22.850 7.480 23.130 7.760 ;
        RECT 38.800 7.480 39.080 7.760 ;
        RECT 53.630 7.480 53.910 7.760 ;
        RECT 22.850 6.820 23.130 7.100 ;
        RECT 38.800 6.820 39.080 7.100 ;
        RECT 53.630 6.820 53.910 7.100 ;
        RECT 26.270 4.770 26.550 5.050 ;
        RECT 26.930 4.770 27.210 5.050 ;
        RECT 27.590 4.770 27.870 5.050 ;
        RECT 32.800 4.740 33.080 5.020 ;
        RECT 33.460 4.740 33.740 5.020 ;
        RECT 34.120 4.740 34.400 5.020 ;
        RECT 36.180 4.740 36.460 5.020 ;
        RECT 42.220 4.770 42.500 5.050 ;
        RECT 42.880 4.770 43.160 5.050 ;
        RECT 43.540 4.770 43.820 5.050 ;
        RECT 48.750 4.740 49.030 5.020 ;
        RECT 49.410 4.740 49.690 5.020 ;
        RECT 50.070 4.740 50.350 5.020 ;
        RECT 57.050 4.770 57.330 5.050 ;
        RECT 57.710 4.770 57.990 5.050 ;
        RECT 58.370 4.770 58.650 5.050 ;
        RECT 63.580 4.740 63.860 5.020 ;
        RECT 64.240 4.740 64.520 5.020 ;
        RECT 64.900 4.740 65.180 5.020 ;
        RECT 66.940 4.740 67.220 5.020 ;
        RECT 67.600 4.740 67.880 5.020 ;
        RECT 68.260 4.740 68.540 5.020 ;
        RECT 4.220 3.470 4.500 3.750 ;
        RECT 4.630 2.810 4.910 3.090 ;
        RECT 22.410 3.470 22.690 3.750 ;
        RECT 22.820 2.810 23.100 3.090 ;
        RECT 38.360 3.470 38.640 3.750 ;
        RECT 38.770 2.810 39.050 3.090 ;
        RECT 96.245 58.795 96.525 59.075 ;
        RECT 96.245 58.135 96.525 58.415 ;
        RECT 96.245 57.475 96.525 57.755 ;
        RECT 96.245 56.815 96.525 57.095 ;
        RECT 96.245 56.155 96.525 56.435 ;
        RECT 96.245 55.495 96.525 55.775 ;
        RECT 96.245 54.835 96.525 55.115 ;
        RECT 96.245 54.175 96.525 54.455 ;
        RECT 96.245 53.515 96.525 53.795 ;
        RECT 96.245 52.855 96.525 53.135 ;
        RECT 96.245 52.195 96.525 52.475 ;
        RECT 96.245 51.535 96.525 51.815 ;
        RECT 96.245 50.875 96.525 51.155 ;
        RECT 96.245 50.215 96.525 50.495 ;
        RECT 106.530 58.795 106.810 59.075 ;
        RECT 106.530 58.135 106.810 58.415 ;
        RECT 106.530 57.475 106.810 57.755 ;
        RECT 106.530 56.815 106.810 57.095 ;
        RECT 106.530 56.155 106.810 56.435 ;
        RECT 106.530 55.495 106.810 55.775 ;
        RECT 106.530 54.835 106.810 55.115 ;
        RECT 106.530 54.175 106.810 54.455 ;
        RECT 106.530 53.515 106.810 53.795 ;
        RECT 106.530 52.855 106.810 53.135 ;
        RECT 106.530 52.195 106.810 52.475 ;
        RECT 106.530 51.535 106.810 51.815 ;
        RECT 106.530 50.875 106.810 51.155 ;
        RECT 106.530 50.215 106.810 50.495 ;
        RECT 100.740 45.155 101.020 45.435 ;
        RECT 101.400 45.155 101.680 45.435 ;
        RECT 102.060 45.155 102.340 45.435 ;
        RECT 100.740 44.495 101.020 44.775 ;
        RECT 101.400 44.495 101.680 44.775 ;
        RECT 102.060 44.495 102.340 44.775 ;
        RECT 100.740 43.835 101.020 44.115 ;
        RECT 101.400 43.835 101.680 44.115 ;
        RECT 102.060 43.835 102.340 44.115 ;
        RECT 111.015 42.455 111.295 42.735 ;
        RECT 111.675 42.455 111.955 42.735 ;
        RECT 112.335 42.455 112.615 42.735 ;
        RECT 111.015 41.795 111.295 42.075 ;
        RECT 111.675 41.795 111.955 42.075 ;
        RECT 112.335 41.795 112.615 42.075 ;
        RECT 111.015 41.135 111.295 41.415 ;
        RECT 111.675 41.135 111.955 41.415 ;
        RECT 112.335 41.135 112.615 41.415 ;
        RECT 111.015 27.655 111.295 27.935 ;
        RECT 111.675 27.655 111.955 27.935 ;
        RECT 112.335 27.655 112.615 27.935 ;
        RECT 111.015 26.995 111.295 27.275 ;
        RECT 111.675 26.995 111.955 27.275 ;
        RECT 112.335 26.995 112.615 27.275 ;
        RECT 111.015 26.335 111.295 26.615 ;
        RECT 111.675 26.335 111.955 26.615 ;
        RECT 112.335 26.335 112.615 26.615 ;
        RECT 100.740 24.955 101.020 25.235 ;
        RECT 101.400 24.955 101.680 25.235 ;
        RECT 102.060 24.955 102.340 25.235 ;
        RECT 100.740 24.295 101.020 24.575 ;
        RECT 101.400 24.295 101.680 24.575 ;
        RECT 102.060 24.295 102.340 24.575 ;
        RECT 100.740 23.635 101.020 23.915 ;
        RECT 101.400 23.635 101.680 23.915 ;
        RECT 102.060 23.635 102.340 23.915 ;
        RECT 116.820 58.795 117.100 59.075 ;
        RECT 116.820 58.135 117.100 58.415 ;
        RECT 116.820 57.475 117.100 57.755 ;
        RECT 116.820 56.815 117.100 57.095 ;
        RECT 116.820 56.155 117.100 56.435 ;
        RECT 116.820 55.495 117.100 55.775 ;
        RECT 116.820 54.835 117.100 55.115 ;
        RECT 116.820 54.175 117.100 54.455 ;
        RECT 116.820 53.515 117.100 53.795 ;
        RECT 116.820 52.855 117.100 53.135 ;
        RECT 116.820 52.195 117.100 52.475 ;
        RECT 116.820 51.535 117.100 51.815 ;
        RECT 116.820 50.875 117.100 51.155 ;
        RECT 116.820 50.215 117.100 50.495 ;
        RECT 127.105 58.795 127.385 59.075 ;
        RECT 128.525 58.795 128.805 59.075 ;
        RECT 127.105 58.135 127.385 58.415 ;
        RECT 128.525 58.135 128.805 58.415 ;
        RECT 127.105 57.475 127.385 57.755 ;
        RECT 128.525 57.475 128.805 57.755 ;
        RECT 127.105 56.815 127.385 57.095 ;
        RECT 128.525 56.815 128.805 57.095 ;
        RECT 127.105 56.155 127.385 56.435 ;
        RECT 128.525 56.155 128.805 56.435 ;
        RECT 127.105 55.495 127.385 55.775 ;
        RECT 128.525 55.495 128.805 55.775 ;
        RECT 127.105 54.835 127.385 55.115 ;
        RECT 128.525 54.835 128.805 55.115 ;
        RECT 127.105 54.175 127.385 54.455 ;
        RECT 128.525 54.175 128.805 54.455 ;
        RECT 127.105 53.515 127.385 53.795 ;
        RECT 128.525 53.515 128.805 53.795 ;
        RECT 127.105 52.855 127.385 53.135 ;
        RECT 128.525 52.855 128.805 53.135 ;
        RECT 127.105 52.195 127.385 52.475 ;
        RECT 128.525 52.195 128.805 52.475 ;
        RECT 127.105 51.535 127.385 51.815 ;
        RECT 128.525 51.535 128.805 51.815 ;
        RECT 127.105 50.875 127.385 51.155 ;
        RECT 128.525 50.875 128.805 51.155 ;
        RECT 127.105 50.215 127.385 50.495 ;
        RECT 128.525 50.215 128.805 50.495 ;
        RECT 133.010 47.855 133.290 48.135 ;
        RECT 133.670 47.855 133.950 48.135 ;
        RECT 134.330 47.855 134.610 48.135 ;
        RECT 133.010 47.195 133.290 47.475 ;
        RECT 133.670 47.195 133.950 47.475 ;
        RECT 134.330 47.195 134.610 47.475 ;
        RECT 133.010 46.535 133.290 46.815 ;
        RECT 133.670 46.535 133.950 46.815 ;
        RECT 134.330 46.535 134.610 46.815 ;
        RECT 121.315 39.755 121.595 40.035 ;
        RECT 121.975 39.755 122.255 40.035 ;
        RECT 122.635 39.755 122.915 40.035 ;
        RECT 121.315 39.095 121.595 39.375 ;
        RECT 121.975 39.095 122.255 39.375 ;
        RECT 122.635 39.095 122.915 39.375 ;
        RECT 121.315 38.435 121.595 38.715 ;
        RECT 121.975 38.435 122.255 38.715 ;
        RECT 122.635 38.435 122.915 38.715 ;
        RECT 121.315 30.355 121.595 30.635 ;
        RECT 121.975 30.355 122.255 30.635 ;
        RECT 122.635 30.355 122.915 30.635 ;
        RECT 121.315 29.695 121.595 29.975 ;
        RECT 121.975 29.695 122.255 29.975 ;
        RECT 122.635 29.695 122.915 29.975 ;
        RECT 121.315 29.035 121.595 29.315 ;
        RECT 121.975 29.035 122.255 29.315 ;
        RECT 122.635 29.035 122.915 29.315 ;
        RECT 133.010 22.255 133.290 22.535 ;
        RECT 133.670 22.255 133.950 22.535 ;
        RECT 134.330 22.255 134.610 22.535 ;
        RECT 133.010 21.595 133.290 21.875 ;
        RECT 133.670 21.595 133.950 21.875 ;
        RECT 134.330 21.595 134.610 21.875 ;
        RECT 133.010 20.935 133.290 21.215 ;
        RECT 133.670 20.935 133.950 21.215 ;
        RECT 134.330 20.935 134.610 21.215 ;
        RECT 72.940 8.140 73.220 8.420 ;
        RECT 87.770 8.140 88.050 8.420 ;
        RECT 72.940 7.480 73.220 7.760 ;
        RECT 87.770 7.480 88.050 7.760 ;
        RECT 72.940 6.820 73.220 7.100 ;
        RECT 87.770 6.820 88.050 7.100 ;
        RECT 70.320 4.740 70.600 5.020 ;
        RECT 76.360 4.770 76.640 5.050 ;
        RECT 77.020 4.770 77.300 5.050 ;
        RECT 77.680 4.770 77.960 5.050 ;
        RECT 82.890 4.740 83.170 5.020 ;
        RECT 83.550 4.740 83.830 5.020 ;
        RECT 84.210 4.740 84.490 5.020 ;
        RECT 91.190 4.770 91.470 5.050 ;
        RECT 91.850 4.770 92.130 5.050 ;
        RECT 92.510 4.770 92.790 5.050 ;
        RECT 97.720 4.740 98.000 5.020 ;
        RECT 98.380 4.740 98.660 5.020 ;
        RECT 99.040 4.740 99.320 5.020 ;
        RECT 101.080 4.740 101.360 5.020 ;
        RECT 101.740 4.740 102.020 5.020 ;
        RECT 102.400 4.740 102.680 5.020 ;
        RECT 53.190 3.470 53.470 3.750 ;
        RECT 53.600 2.810 53.880 3.090 ;
        RECT 72.500 3.470 72.780 3.750 ;
        RECT 72.910 2.810 73.190 3.090 ;
        RECT 138.815 58.795 139.095 59.075 ;
        RECT 138.815 58.135 139.095 58.415 ;
        RECT 138.815 57.475 139.095 57.755 ;
        RECT 138.815 56.815 139.095 57.095 ;
        RECT 138.815 56.155 139.095 56.435 ;
        RECT 138.815 55.495 139.095 55.775 ;
        RECT 138.815 54.835 139.095 55.115 ;
        RECT 138.815 54.175 139.095 54.455 ;
        RECT 138.815 53.515 139.095 53.795 ;
        RECT 138.815 52.855 139.095 53.135 ;
        RECT 138.815 52.195 139.095 52.475 ;
        RECT 138.815 51.535 139.095 51.815 ;
        RECT 138.815 50.875 139.095 51.155 ;
        RECT 138.815 50.215 139.095 50.495 ;
        RECT 149.100 58.795 149.380 59.075 ;
        RECT 149.100 58.135 149.380 58.415 ;
        RECT 149.100 57.475 149.380 57.755 ;
        RECT 149.100 56.815 149.380 57.095 ;
        RECT 149.100 56.155 149.380 56.435 ;
        RECT 149.100 55.495 149.380 55.775 ;
        RECT 149.100 54.835 149.380 55.115 ;
        RECT 149.100 54.175 149.380 54.455 ;
        RECT 149.100 53.515 149.380 53.795 ;
        RECT 149.100 52.855 149.380 53.135 ;
        RECT 149.100 52.195 149.380 52.475 ;
        RECT 149.100 51.535 149.380 51.815 ;
        RECT 149.100 50.875 149.380 51.155 ;
        RECT 149.100 50.215 149.380 50.495 ;
        RECT 143.310 45.155 143.590 45.435 ;
        RECT 143.970 45.155 144.250 45.435 ;
        RECT 144.630 45.155 144.910 45.435 ;
        RECT 143.310 44.495 143.590 44.775 ;
        RECT 143.970 44.495 144.250 44.775 ;
        RECT 144.630 44.495 144.910 44.775 ;
        RECT 143.310 43.835 143.590 44.115 ;
        RECT 143.970 43.835 144.250 44.115 ;
        RECT 144.630 43.835 144.910 44.115 ;
        RECT 153.585 42.455 153.865 42.735 ;
        RECT 154.245 42.455 154.525 42.735 ;
        RECT 154.905 42.455 155.185 42.735 ;
        RECT 153.585 41.795 153.865 42.075 ;
        RECT 154.245 41.795 154.525 42.075 ;
        RECT 154.905 41.795 155.185 42.075 ;
        RECT 153.585 41.135 153.865 41.415 ;
        RECT 154.245 41.135 154.525 41.415 ;
        RECT 154.905 41.135 155.185 41.415 ;
        RECT 153.585 27.655 153.865 27.935 ;
        RECT 154.245 27.655 154.525 27.935 ;
        RECT 154.905 27.655 155.185 27.935 ;
        RECT 153.585 26.995 153.865 27.275 ;
        RECT 154.245 26.995 154.525 27.275 ;
        RECT 154.905 26.995 155.185 27.275 ;
        RECT 153.585 26.335 153.865 26.615 ;
        RECT 154.245 26.335 154.525 26.615 ;
        RECT 154.905 26.335 155.185 26.615 ;
        RECT 143.310 24.955 143.590 25.235 ;
        RECT 143.970 24.955 144.250 25.235 ;
        RECT 144.630 24.955 144.910 25.235 ;
        RECT 143.310 24.295 143.590 24.575 ;
        RECT 143.970 24.295 144.250 24.575 ;
        RECT 144.630 24.295 144.910 24.575 ;
        RECT 143.310 23.635 143.590 23.915 ;
        RECT 143.970 23.635 144.250 23.915 ;
        RECT 144.630 23.635 144.910 23.915 ;
        RECT 159.390 58.795 159.670 59.075 ;
        RECT 159.390 58.135 159.670 58.415 ;
        RECT 159.390 57.475 159.670 57.755 ;
        RECT 159.390 56.815 159.670 57.095 ;
        RECT 159.390 56.155 159.670 56.435 ;
        RECT 159.390 55.495 159.670 55.775 ;
        RECT 159.390 54.835 159.670 55.115 ;
        RECT 159.390 54.175 159.670 54.455 ;
        RECT 159.390 53.515 159.670 53.795 ;
        RECT 159.390 52.855 159.670 53.135 ;
        RECT 159.390 52.195 159.670 52.475 ;
        RECT 159.390 51.535 159.670 51.815 ;
        RECT 159.390 50.875 159.670 51.155 ;
        RECT 159.390 50.215 159.670 50.495 ;
        RECT 169.675 58.795 169.955 59.075 ;
        RECT 171.095 58.795 171.375 59.075 ;
        RECT 169.675 58.135 169.955 58.415 ;
        RECT 171.095 58.135 171.375 58.415 ;
        RECT 169.675 57.475 169.955 57.755 ;
        RECT 171.095 57.475 171.375 57.755 ;
        RECT 169.675 56.815 169.955 57.095 ;
        RECT 171.095 56.815 171.375 57.095 ;
        RECT 169.675 56.155 169.955 56.435 ;
        RECT 171.095 56.155 171.375 56.435 ;
        RECT 169.675 55.495 169.955 55.775 ;
        RECT 171.095 55.495 171.375 55.775 ;
        RECT 169.675 54.835 169.955 55.115 ;
        RECT 171.095 54.835 171.375 55.115 ;
        RECT 169.675 54.175 169.955 54.455 ;
        RECT 171.095 54.175 171.375 54.455 ;
        RECT 169.675 53.515 169.955 53.795 ;
        RECT 171.095 53.515 171.375 53.795 ;
        RECT 169.675 52.855 169.955 53.135 ;
        RECT 171.095 52.855 171.375 53.135 ;
        RECT 169.675 52.195 169.955 52.475 ;
        RECT 171.095 52.195 171.375 52.475 ;
        RECT 169.675 51.535 169.955 51.815 ;
        RECT 171.095 51.535 171.375 51.815 ;
        RECT 169.675 50.875 169.955 51.155 ;
        RECT 171.095 50.875 171.375 51.155 ;
        RECT 169.675 50.215 169.955 50.495 ;
        RECT 171.095 50.215 171.375 50.495 ;
        RECT 175.580 47.855 175.860 48.135 ;
        RECT 176.240 47.855 176.520 48.135 ;
        RECT 176.900 47.855 177.180 48.135 ;
        RECT 175.580 47.195 175.860 47.475 ;
        RECT 176.240 47.195 176.520 47.475 ;
        RECT 176.900 47.195 177.180 47.475 ;
        RECT 175.580 46.535 175.860 46.815 ;
        RECT 176.240 46.535 176.520 46.815 ;
        RECT 176.900 46.535 177.180 46.815 ;
        RECT 163.885 39.755 164.165 40.035 ;
        RECT 164.545 39.755 164.825 40.035 ;
        RECT 165.205 39.755 165.485 40.035 ;
        RECT 163.885 39.095 164.165 39.375 ;
        RECT 164.545 39.095 164.825 39.375 ;
        RECT 165.205 39.095 165.485 39.375 ;
        RECT 163.885 38.435 164.165 38.715 ;
        RECT 164.545 38.435 164.825 38.715 ;
        RECT 165.205 38.435 165.485 38.715 ;
        RECT 163.885 30.355 164.165 30.635 ;
        RECT 164.545 30.355 164.825 30.635 ;
        RECT 165.205 30.355 165.485 30.635 ;
        RECT 163.885 29.695 164.165 29.975 ;
        RECT 164.545 29.695 164.825 29.975 ;
        RECT 165.205 29.695 165.485 29.975 ;
        RECT 163.885 29.035 164.165 29.315 ;
        RECT 164.545 29.035 164.825 29.315 ;
        RECT 165.205 29.035 165.485 29.315 ;
        RECT 175.580 22.255 175.860 22.535 ;
        RECT 176.240 22.255 176.520 22.535 ;
        RECT 176.900 22.255 177.180 22.535 ;
        RECT 175.580 21.595 175.860 21.875 ;
        RECT 176.240 21.595 176.520 21.875 ;
        RECT 176.900 21.595 177.180 21.875 ;
        RECT 175.580 20.935 175.860 21.215 ;
        RECT 176.240 20.935 176.520 21.215 ;
        RECT 176.900 20.935 177.180 21.215 ;
        RECT 107.080 8.140 107.360 8.420 ;
        RECT 121.910 8.140 122.190 8.420 ;
        RECT 107.080 7.480 107.360 7.760 ;
        RECT 121.910 7.480 122.190 7.760 ;
        RECT 107.080 6.820 107.360 7.100 ;
        RECT 121.910 6.820 122.190 7.100 ;
        RECT 104.460 4.740 104.740 5.020 ;
        RECT 110.500 4.770 110.780 5.050 ;
        RECT 111.160 4.770 111.440 5.050 ;
        RECT 111.820 4.770 112.100 5.050 ;
        RECT 117.030 4.740 117.310 5.020 ;
        RECT 117.690 4.740 117.970 5.020 ;
        RECT 118.350 4.740 118.630 5.020 ;
        RECT 125.330 4.770 125.610 5.050 ;
        RECT 125.990 4.770 126.270 5.050 ;
        RECT 126.650 4.770 126.930 5.050 ;
        RECT 131.860 4.740 132.140 5.020 ;
        RECT 132.520 4.740 132.800 5.020 ;
        RECT 133.180 4.740 133.460 5.020 ;
        RECT 135.240 4.740 135.520 5.020 ;
        RECT 136.240 4.740 136.520 5.020 ;
        RECT 136.900 4.740 137.180 5.020 ;
        RECT 137.560 4.740 137.840 5.020 ;
        RECT 138.480 4.740 138.760 5.020 ;
        RECT 139.140 4.740 139.420 5.020 ;
        RECT 139.800 4.740 140.080 5.020 ;
        RECT 140.820 4.740 141.100 5.020 ;
        RECT 141.480 4.740 141.760 5.020 ;
        RECT 142.140 4.740 142.420 5.020 ;
        RECT 87.330 3.470 87.610 3.750 ;
        RECT 87.740 2.810 88.020 3.090 ;
        RECT 106.640 3.470 106.920 3.750 ;
        RECT 107.050 2.810 107.330 3.090 ;
        RECT 181.385 58.795 181.665 59.075 ;
        RECT 181.385 58.135 181.665 58.415 ;
        RECT 181.385 57.475 181.665 57.755 ;
        RECT 181.385 56.815 181.665 57.095 ;
        RECT 181.385 56.155 181.665 56.435 ;
        RECT 181.385 55.495 181.665 55.775 ;
        RECT 181.385 54.835 181.665 55.115 ;
        RECT 181.385 54.175 181.665 54.455 ;
        RECT 181.385 53.515 181.665 53.795 ;
        RECT 181.385 52.855 181.665 53.135 ;
        RECT 181.385 52.195 181.665 52.475 ;
        RECT 181.385 51.535 181.665 51.815 ;
        RECT 181.385 50.875 181.665 51.155 ;
        RECT 181.385 50.215 181.665 50.495 ;
        RECT 191.670 58.795 191.950 59.075 ;
        RECT 191.670 58.135 191.950 58.415 ;
        RECT 191.670 57.475 191.950 57.755 ;
        RECT 191.670 56.815 191.950 57.095 ;
        RECT 191.670 56.155 191.950 56.435 ;
        RECT 191.670 55.495 191.950 55.775 ;
        RECT 191.670 54.835 191.950 55.115 ;
        RECT 191.670 54.175 191.950 54.455 ;
        RECT 191.670 53.515 191.950 53.795 ;
        RECT 191.670 52.855 191.950 53.135 ;
        RECT 191.670 52.195 191.950 52.475 ;
        RECT 191.670 51.535 191.950 51.815 ;
        RECT 191.670 50.875 191.950 51.155 ;
        RECT 191.670 50.215 191.950 50.495 ;
        RECT 185.880 45.155 186.160 45.435 ;
        RECT 186.540 45.155 186.820 45.435 ;
        RECT 187.200 45.155 187.480 45.435 ;
        RECT 185.880 44.495 186.160 44.775 ;
        RECT 186.540 44.495 186.820 44.775 ;
        RECT 187.200 44.495 187.480 44.775 ;
        RECT 185.880 43.835 186.160 44.115 ;
        RECT 186.540 43.835 186.820 44.115 ;
        RECT 187.200 43.835 187.480 44.115 ;
        RECT 196.155 42.455 196.435 42.735 ;
        RECT 196.815 42.455 197.095 42.735 ;
        RECT 197.475 42.455 197.755 42.735 ;
        RECT 196.155 41.795 196.435 42.075 ;
        RECT 196.815 41.795 197.095 42.075 ;
        RECT 197.475 41.795 197.755 42.075 ;
        RECT 196.155 41.135 196.435 41.415 ;
        RECT 196.815 41.135 197.095 41.415 ;
        RECT 197.475 41.135 197.755 41.415 ;
        RECT 196.155 27.655 196.435 27.935 ;
        RECT 196.815 27.655 197.095 27.935 ;
        RECT 197.475 27.655 197.755 27.935 ;
        RECT 196.155 26.995 196.435 27.275 ;
        RECT 196.815 26.995 197.095 27.275 ;
        RECT 197.475 26.995 197.755 27.275 ;
        RECT 196.155 26.335 196.435 26.615 ;
        RECT 196.815 26.335 197.095 26.615 ;
        RECT 197.475 26.335 197.755 26.615 ;
        RECT 185.880 24.955 186.160 25.235 ;
        RECT 186.540 24.955 186.820 25.235 ;
        RECT 187.200 24.955 187.480 25.235 ;
        RECT 185.880 24.295 186.160 24.575 ;
        RECT 186.540 24.295 186.820 24.575 ;
        RECT 187.200 24.295 187.480 24.575 ;
        RECT 185.880 23.635 186.160 23.915 ;
        RECT 186.540 23.635 186.820 23.915 ;
        RECT 187.200 23.635 187.480 23.915 ;
        RECT 201.960 58.795 202.240 59.075 ;
        RECT 201.960 58.135 202.240 58.415 ;
        RECT 201.960 57.475 202.240 57.755 ;
        RECT 201.960 56.815 202.240 57.095 ;
        RECT 201.960 56.155 202.240 56.435 ;
        RECT 201.960 55.495 202.240 55.775 ;
        RECT 201.960 54.835 202.240 55.115 ;
        RECT 201.960 54.175 202.240 54.455 ;
        RECT 201.960 53.515 202.240 53.795 ;
        RECT 201.960 52.855 202.240 53.135 ;
        RECT 201.960 52.195 202.240 52.475 ;
        RECT 201.960 51.535 202.240 51.815 ;
        RECT 201.960 50.875 202.240 51.155 ;
        RECT 201.960 50.215 202.240 50.495 ;
        RECT 212.245 58.795 212.525 59.075 ;
        RECT 213.665 58.795 213.945 59.075 ;
        RECT 212.245 58.135 212.525 58.415 ;
        RECT 213.665 58.135 213.945 58.415 ;
        RECT 212.245 57.475 212.525 57.755 ;
        RECT 213.665 57.475 213.945 57.755 ;
        RECT 212.245 56.815 212.525 57.095 ;
        RECT 213.665 56.815 213.945 57.095 ;
        RECT 212.245 56.155 212.525 56.435 ;
        RECT 213.665 56.155 213.945 56.435 ;
        RECT 212.245 55.495 212.525 55.775 ;
        RECT 213.665 55.495 213.945 55.775 ;
        RECT 212.245 54.835 212.525 55.115 ;
        RECT 213.665 54.835 213.945 55.115 ;
        RECT 212.245 54.175 212.525 54.455 ;
        RECT 213.665 54.175 213.945 54.455 ;
        RECT 212.245 53.515 212.525 53.795 ;
        RECT 213.665 53.515 213.945 53.795 ;
        RECT 212.245 52.855 212.525 53.135 ;
        RECT 213.665 52.855 213.945 53.135 ;
        RECT 212.245 52.195 212.525 52.475 ;
        RECT 213.665 52.195 213.945 52.475 ;
        RECT 212.245 51.535 212.525 51.815 ;
        RECT 213.665 51.535 213.945 51.815 ;
        RECT 212.245 50.875 212.525 51.155 ;
        RECT 213.665 50.875 213.945 51.155 ;
        RECT 212.245 50.215 212.525 50.495 ;
        RECT 213.665 50.215 213.945 50.495 ;
        RECT 218.150 47.855 218.430 48.135 ;
        RECT 218.810 47.855 219.090 48.135 ;
        RECT 219.470 47.855 219.750 48.135 ;
        RECT 218.150 47.195 218.430 47.475 ;
        RECT 218.810 47.195 219.090 47.475 ;
        RECT 219.470 47.195 219.750 47.475 ;
        RECT 218.150 46.535 218.430 46.815 ;
        RECT 218.810 46.535 219.090 46.815 ;
        RECT 219.470 46.535 219.750 46.815 ;
        RECT 206.455 39.755 206.735 40.035 ;
        RECT 207.115 39.755 207.395 40.035 ;
        RECT 207.775 39.755 208.055 40.035 ;
        RECT 206.455 39.095 206.735 39.375 ;
        RECT 207.115 39.095 207.395 39.375 ;
        RECT 207.775 39.095 208.055 39.375 ;
        RECT 206.455 38.435 206.735 38.715 ;
        RECT 207.115 38.435 207.395 38.715 ;
        RECT 207.775 38.435 208.055 38.715 ;
        RECT 206.455 30.355 206.735 30.635 ;
        RECT 207.115 30.355 207.395 30.635 ;
        RECT 207.775 30.355 208.055 30.635 ;
        RECT 206.455 29.695 206.735 29.975 ;
        RECT 207.115 29.695 207.395 29.975 ;
        RECT 207.775 29.695 208.055 29.975 ;
        RECT 206.455 29.035 206.735 29.315 ;
        RECT 207.115 29.035 207.395 29.315 ;
        RECT 207.775 29.035 208.055 29.315 ;
        RECT 218.150 22.255 218.430 22.535 ;
        RECT 218.810 22.255 219.090 22.535 ;
        RECT 219.470 22.255 219.750 22.535 ;
        RECT 218.150 21.595 218.430 21.875 ;
        RECT 218.810 21.595 219.090 21.875 ;
        RECT 219.470 21.595 219.750 21.875 ;
        RECT 218.150 20.935 218.430 21.215 ;
        RECT 218.810 20.935 219.090 21.215 ;
        RECT 219.470 20.935 219.750 21.215 ;
        RECT 144.080 4.740 144.360 5.020 ;
        RECT 144.740 4.740 145.020 5.020 ;
        RECT 145.400 4.740 145.680 5.020 ;
        RECT 146.320 4.740 146.600 5.020 ;
        RECT 146.980 4.740 147.260 5.020 ;
        RECT 147.640 4.740 147.920 5.020 ;
        RECT 148.560 4.740 148.840 5.020 ;
        RECT 149.220 4.740 149.500 5.020 ;
        RECT 149.880 4.740 150.160 5.020 ;
        RECT 150.800 4.740 151.080 5.020 ;
        RECT 151.460 4.740 151.740 5.020 ;
        RECT 152.120 4.740 152.400 5.020 ;
        RECT 153.040 4.740 153.320 5.020 ;
        RECT 153.700 4.740 153.980 5.020 ;
        RECT 154.360 4.740 154.640 5.020 ;
        RECT 155.400 4.740 155.680 5.020 ;
        RECT 156.400 4.740 156.680 5.020 ;
        RECT 157.060 4.740 157.340 5.020 ;
        RECT 157.720 4.740 158.000 5.020 ;
        RECT 158.640 4.740 158.920 5.020 ;
        RECT 159.300 4.740 159.580 5.020 ;
        RECT 159.960 4.740 160.240 5.020 ;
        RECT 160.880 4.740 161.160 5.020 ;
        RECT 161.540 4.740 161.820 5.020 ;
        RECT 162.200 4.740 162.480 5.020 ;
        RECT 163.120 4.740 163.400 5.020 ;
        RECT 163.780 4.740 164.060 5.020 ;
        RECT 164.440 4.740 164.720 5.020 ;
        RECT 165.360 4.740 165.640 5.020 ;
        RECT 166.020 4.740 166.300 5.020 ;
        RECT 166.680 4.740 166.960 5.020 ;
        RECT 167.600 4.740 167.880 5.020 ;
        RECT 168.260 4.740 168.540 5.020 ;
        RECT 168.920 4.740 169.200 5.020 ;
        RECT 169.840 4.740 170.120 5.020 ;
        RECT 170.500 4.740 170.780 5.020 ;
        RECT 171.160 4.740 171.440 5.020 ;
        RECT 172.080 4.740 172.360 5.020 ;
        RECT 172.740 4.740 173.020 5.020 ;
        RECT 173.400 4.740 173.680 5.020 ;
        RECT 174.320 4.740 174.600 5.020 ;
        RECT 174.980 4.740 175.260 5.020 ;
        RECT 175.640 4.740 175.920 5.020 ;
        RECT 176.680 4.740 176.960 5.020 ;
        RECT 177.680 4.740 177.960 5.020 ;
        RECT 178.340 4.740 178.620 5.020 ;
        RECT 179.000 4.740 179.280 5.020 ;
        RECT 179.920 4.740 180.200 5.020 ;
        RECT 180.580 4.740 180.860 5.020 ;
        RECT 181.240 4.740 181.520 5.020 ;
        RECT 182.260 4.740 182.540 5.020 ;
        RECT 182.920 4.740 183.200 5.020 ;
        RECT 183.580 4.740 183.860 5.020 ;
        RECT 223.955 58.795 224.235 59.075 ;
        RECT 223.955 58.135 224.235 58.415 ;
        RECT 223.955 57.475 224.235 57.755 ;
        RECT 223.955 56.815 224.235 57.095 ;
        RECT 223.955 56.155 224.235 56.435 ;
        RECT 223.955 55.495 224.235 55.775 ;
        RECT 223.955 54.835 224.235 55.115 ;
        RECT 223.955 54.175 224.235 54.455 ;
        RECT 223.955 53.515 224.235 53.795 ;
        RECT 223.955 52.855 224.235 53.135 ;
        RECT 223.955 52.195 224.235 52.475 ;
        RECT 223.955 51.535 224.235 51.815 ;
        RECT 223.955 50.875 224.235 51.155 ;
        RECT 223.955 50.215 224.235 50.495 ;
        RECT 234.240 58.795 234.520 59.075 ;
        RECT 234.240 58.135 234.520 58.415 ;
        RECT 234.240 57.475 234.520 57.755 ;
        RECT 234.240 56.815 234.520 57.095 ;
        RECT 234.240 56.155 234.520 56.435 ;
        RECT 234.240 55.495 234.520 55.775 ;
        RECT 234.240 54.835 234.520 55.115 ;
        RECT 234.240 54.175 234.520 54.455 ;
        RECT 234.240 53.515 234.520 53.795 ;
        RECT 234.240 52.855 234.520 53.135 ;
        RECT 234.240 52.195 234.520 52.475 ;
        RECT 234.240 51.535 234.520 51.815 ;
        RECT 234.240 50.875 234.520 51.155 ;
        RECT 234.240 50.215 234.520 50.495 ;
        RECT 228.450 45.155 228.730 45.435 ;
        RECT 229.110 45.155 229.390 45.435 ;
        RECT 229.770 45.155 230.050 45.435 ;
        RECT 228.450 44.495 228.730 44.775 ;
        RECT 229.110 44.495 229.390 44.775 ;
        RECT 229.770 44.495 230.050 44.775 ;
        RECT 228.450 43.835 228.730 44.115 ;
        RECT 229.110 43.835 229.390 44.115 ;
        RECT 229.770 43.835 230.050 44.115 ;
        RECT 238.725 42.455 239.005 42.735 ;
        RECT 239.385 42.455 239.665 42.735 ;
        RECT 240.045 42.455 240.325 42.735 ;
        RECT 238.725 41.795 239.005 42.075 ;
        RECT 239.385 41.795 239.665 42.075 ;
        RECT 240.045 41.795 240.325 42.075 ;
        RECT 238.725 41.135 239.005 41.415 ;
        RECT 239.385 41.135 239.665 41.415 ;
        RECT 240.045 41.135 240.325 41.415 ;
        RECT 238.725 27.655 239.005 27.935 ;
        RECT 239.385 27.655 239.665 27.935 ;
        RECT 240.045 27.655 240.325 27.935 ;
        RECT 238.725 26.995 239.005 27.275 ;
        RECT 239.385 26.995 239.665 27.275 ;
        RECT 240.045 26.995 240.325 27.275 ;
        RECT 238.725 26.335 239.005 26.615 ;
        RECT 239.385 26.335 239.665 26.615 ;
        RECT 240.045 26.335 240.325 26.615 ;
        RECT 228.450 24.955 228.730 25.235 ;
        RECT 229.110 24.955 229.390 25.235 ;
        RECT 229.770 24.955 230.050 25.235 ;
        RECT 228.450 24.295 228.730 24.575 ;
        RECT 229.110 24.295 229.390 24.575 ;
        RECT 229.770 24.295 230.050 24.575 ;
        RECT 228.450 23.635 228.730 23.915 ;
        RECT 229.110 23.635 229.390 23.915 ;
        RECT 229.770 23.635 230.050 23.915 ;
        RECT 244.530 58.795 244.810 59.075 ;
        RECT 244.530 58.135 244.810 58.415 ;
        RECT 244.530 57.475 244.810 57.755 ;
        RECT 244.530 56.815 244.810 57.095 ;
        RECT 244.530 56.155 244.810 56.435 ;
        RECT 244.530 55.495 244.810 55.775 ;
        RECT 244.530 54.835 244.810 55.115 ;
        RECT 244.530 54.175 244.810 54.455 ;
        RECT 244.530 53.515 244.810 53.795 ;
        RECT 244.530 52.855 244.810 53.135 ;
        RECT 244.530 52.195 244.810 52.475 ;
        RECT 244.530 51.535 244.810 51.815 ;
        RECT 244.530 50.875 244.810 51.155 ;
        RECT 244.530 50.215 244.810 50.495 ;
        RECT 254.815 58.795 255.095 59.075 ;
        RECT 256.235 58.795 256.515 59.075 ;
        RECT 254.815 58.135 255.095 58.415 ;
        RECT 256.235 58.135 256.515 58.415 ;
        RECT 254.815 57.475 255.095 57.755 ;
        RECT 256.235 57.475 256.515 57.755 ;
        RECT 254.815 56.815 255.095 57.095 ;
        RECT 256.235 56.815 256.515 57.095 ;
        RECT 254.815 56.155 255.095 56.435 ;
        RECT 256.235 56.155 256.515 56.435 ;
        RECT 254.815 55.495 255.095 55.775 ;
        RECT 256.235 55.495 256.515 55.775 ;
        RECT 254.815 54.835 255.095 55.115 ;
        RECT 256.235 54.835 256.515 55.115 ;
        RECT 254.815 54.175 255.095 54.455 ;
        RECT 256.235 54.175 256.515 54.455 ;
        RECT 254.815 53.515 255.095 53.795 ;
        RECT 256.235 53.515 256.515 53.795 ;
        RECT 254.815 52.855 255.095 53.135 ;
        RECT 256.235 52.855 256.515 53.135 ;
        RECT 254.815 52.195 255.095 52.475 ;
        RECT 256.235 52.195 256.515 52.475 ;
        RECT 254.815 51.535 255.095 51.815 ;
        RECT 256.235 51.535 256.515 51.815 ;
        RECT 254.815 50.875 255.095 51.155 ;
        RECT 256.235 50.875 256.515 51.155 ;
        RECT 254.815 50.215 255.095 50.495 ;
        RECT 256.235 50.215 256.515 50.495 ;
        RECT 260.720 47.855 261.000 48.135 ;
        RECT 261.380 47.855 261.660 48.135 ;
        RECT 262.040 47.855 262.320 48.135 ;
        RECT 260.720 47.195 261.000 47.475 ;
        RECT 261.380 47.195 261.660 47.475 ;
        RECT 262.040 47.195 262.320 47.475 ;
        RECT 260.720 46.535 261.000 46.815 ;
        RECT 261.380 46.535 261.660 46.815 ;
        RECT 262.040 46.535 262.320 46.815 ;
        RECT 249.025 39.755 249.305 40.035 ;
        RECT 249.685 39.755 249.965 40.035 ;
        RECT 250.345 39.755 250.625 40.035 ;
        RECT 249.025 39.095 249.305 39.375 ;
        RECT 249.685 39.095 249.965 39.375 ;
        RECT 250.345 39.095 250.625 39.375 ;
        RECT 249.025 38.435 249.305 38.715 ;
        RECT 249.685 38.435 249.965 38.715 ;
        RECT 250.345 38.435 250.625 38.715 ;
        RECT 249.025 30.355 249.305 30.635 ;
        RECT 249.685 30.355 249.965 30.635 ;
        RECT 250.345 30.355 250.625 30.635 ;
        RECT 249.025 29.695 249.305 29.975 ;
        RECT 249.685 29.695 249.965 29.975 ;
        RECT 250.345 29.695 250.625 29.975 ;
        RECT 249.025 29.035 249.305 29.315 ;
        RECT 249.685 29.035 249.965 29.315 ;
        RECT 250.345 29.035 250.625 29.315 ;
        RECT 260.720 22.255 261.000 22.535 ;
        RECT 261.380 22.255 261.660 22.535 ;
        RECT 262.040 22.255 262.320 22.535 ;
        RECT 260.720 21.595 261.000 21.875 ;
        RECT 261.380 21.595 261.660 21.875 ;
        RECT 262.040 21.595 262.320 21.875 ;
        RECT 260.720 20.935 261.000 21.215 ;
        RECT 261.380 20.935 261.660 21.215 ;
        RECT 262.040 20.935 262.320 21.215 ;
        RECT 185.520 4.740 185.800 5.020 ;
        RECT 186.180 4.740 186.460 5.020 ;
        RECT 186.840 4.740 187.120 5.020 ;
        RECT 187.760 4.740 188.040 5.020 ;
        RECT 188.420 4.740 188.700 5.020 ;
        RECT 189.080 4.740 189.360 5.020 ;
        RECT 190.000 4.740 190.280 5.020 ;
        RECT 190.660 4.740 190.940 5.020 ;
        RECT 191.320 4.740 191.600 5.020 ;
        RECT 192.240 4.740 192.520 5.020 ;
        RECT 192.900 4.740 193.180 5.020 ;
        RECT 193.560 4.740 193.840 5.020 ;
        RECT 194.480 4.740 194.760 5.020 ;
        RECT 195.140 4.740 195.420 5.020 ;
        RECT 195.800 4.740 196.080 5.020 ;
        RECT 196.840 4.740 197.120 5.020 ;
        RECT 197.840 4.740 198.120 5.020 ;
        RECT 198.500 4.740 198.780 5.020 ;
        RECT 199.160 4.740 199.440 5.020 ;
        RECT 200.080 4.740 200.360 5.020 ;
        RECT 200.740 4.740 201.020 5.020 ;
        RECT 201.400 4.740 201.680 5.020 ;
        RECT 202.320 4.740 202.600 5.020 ;
        RECT 202.980 4.740 203.260 5.020 ;
        RECT 203.640 4.740 203.920 5.020 ;
        RECT 204.560 4.740 204.840 5.020 ;
        RECT 205.220 4.740 205.500 5.020 ;
        RECT 205.880 4.740 206.160 5.020 ;
        RECT 206.800 4.740 207.080 5.020 ;
        RECT 207.460 4.740 207.740 5.020 ;
        RECT 208.120 4.740 208.400 5.020 ;
        RECT 209.040 4.740 209.320 5.020 ;
        RECT 209.700 4.740 209.980 5.020 ;
        RECT 210.360 4.740 210.640 5.020 ;
        RECT 211.280 4.740 211.560 5.020 ;
        RECT 211.940 4.740 212.220 5.020 ;
        RECT 212.600 4.740 212.880 5.020 ;
        RECT 213.520 4.740 213.800 5.020 ;
        RECT 214.180 4.740 214.460 5.020 ;
        RECT 214.840 4.740 215.120 5.020 ;
        RECT 215.760 4.740 216.040 5.020 ;
        RECT 216.420 4.740 216.700 5.020 ;
        RECT 217.080 4.740 217.360 5.020 ;
        RECT 218.120 4.740 218.400 5.020 ;
        RECT 219.120 4.740 219.400 5.020 ;
        RECT 219.780 4.740 220.060 5.020 ;
        RECT 220.440 4.740 220.720 5.020 ;
        RECT 221.360 4.740 221.640 5.020 ;
        RECT 222.020 4.740 222.300 5.020 ;
        RECT 222.680 4.740 222.960 5.020 ;
        RECT 223.600 4.740 223.880 5.020 ;
        RECT 224.260 4.740 224.540 5.020 ;
        RECT 224.920 4.740 225.200 5.020 ;
        RECT 225.940 4.740 226.220 5.020 ;
        RECT 226.600 4.740 226.880 5.020 ;
        RECT 227.260 4.740 227.540 5.020 ;
        RECT 266.525 58.795 266.805 59.075 ;
        RECT 266.525 58.135 266.805 58.415 ;
        RECT 266.525 57.475 266.805 57.755 ;
        RECT 266.525 56.815 266.805 57.095 ;
        RECT 266.525 56.155 266.805 56.435 ;
        RECT 266.525 55.495 266.805 55.775 ;
        RECT 266.525 54.835 266.805 55.115 ;
        RECT 266.525 54.175 266.805 54.455 ;
        RECT 266.525 53.515 266.805 53.795 ;
        RECT 266.525 52.855 266.805 53.135 ;
        RECT 266.525 52.195 266.805 52.475 ;
        RECT 266.525 51.535 266.805 51.815 ;
        RECT 266.525 50.875 266.805 51.155 ;
        RECT 266.525 50.215 266.805 50.495 ;
        RECT 276.810 58.795 277.090 59.075 ;
        RECT 276.810 58.135 277.090 58.415 ;
        RECT 276.810 57.475 277.090 57.755 ;
        RECT 276.810 56.815 277.090 57.095 ;
        RECT 276.810 56.155 277.090 56.435 ;
        RECT 276.810 55.495 277.090 55.775 ;
        RECT 276.810 54.835 277.090 55.115 ;
        RECT 276.810 54.175 277.090 54.455 ;
        RECT 276.810 53.515 277.090 53.795 ;
        RECT 276.810 52.855 277.090 53.135 ;
        RECT 276.810 52.195 277.090 52.475 ;
        RECT 276.810 51.535 277.090 51.815 ;
        RECT 276.810 50.875 277.090 51.155 ;
        RECT 276.810 50.215 277.090 50.495 ;
        RECT 271.020 45.155 271.300 45.435 ;
        RECT 271.680 45.155 271.960 45.435 ;
        RECT 272.340 45.155 272.620 45.435 ;
        RECT 271.020 44.495 271.300 44.775 ;
        RECT 271.680 44.495 271.960 44.775 ;
        RECT 272.340 44.495 272.620 44.775 ;
        RECT 271.020 43.835 271.300 44.115 ;
        RECT 271.680 43.835 271.960 44.115 ;
        RECT 272.340 43.835 272.620 44.115 ;
        RECT 281.295 42.455 281.575 42.735 ;
        RECT 281.955 42.455 282.235 42.735 ;
        RECT 282.615 42.455 282.895 42.735 ;
        RECT 281.295 41.795 281.575 42.075 ;
        RECT 281.955 41.795 282.235 42.075 ;
        RECT 282.615 41.795 282.895 42.075 ;
        RECT 281.295 41.135 281.575 41.415 ;
        RECT 281.955 41.135 282.235 41.415 ;
        RECT 282.615 41.135 282.895 41.415 ;
        RECT 281.295 27.655 281.575 27.935 ;
        RECT 281.955 27.655 282.235 27.935 ;
        RECT 282.615 27.655 282.895 27.935 ;
        RECT 281.295 26.995 281.575 27.275 ;
        RECT 281.955 26.995 282.235 27.275 ;
        RECT 282.615 26.995 282.895 27.275 ;
        RECT 281.295 26.335 281.575 26.615 ;
        RECT 281.955 26.335 282.235 26.615 ;
        RECT 282.615 26.335 282.895 26.615 ;
        RECT 271.020 24.955 271.300 25.235 ;
        RECT 271.680 24.955 271.960 25.235 ;
        RECT 272.340 24.955 272.620 25.235 ;
        RECT 271.020 24.295 271.300 24.575 ;
        RECT 271.680 24.295 271.960 24.575 ;
        RECT 272.340 24.295 272.620 24.575 ;
        RECT 271.020 23.635 271.300 23.915 ;
        RECT 271.680 23.635 271.960 23.915 ;
        RECT 272.340 23.635 272.620 23.915 ;
        RECT 287.100 58.795 287.380 59.075 ;
        RECT 287.100 58.135 287.380 58.415 ;
        RECT 287.100 57.475 287.380 57.755 ;
        RECT 287.100 56.815 287.380 57.095 ;
        RECT 287.100 56.155 287.380 56.435 ;
        RECT 287.100 55.495 287.380 55.775 ;
        RECT 287.100 54.835 287.380 55.115 ;
        RECT 287.100 54.175 287.380 54.455 ;
        RECT 287.100 53.515 287.380 53.795 ;
        RECT 287.100 52.855 287.380 53.135 ;
        RECT 287.100 52.195 287.380 52.475 ;
        RECT 287.100 51.535 287.380 51.815 ;
        RECT 287.100 50.875 287.380 51.155 ;
        RECT 287.100 50.215 287.380 50.495 ;
        RECT 297.385 58.795 297.665 59.075 ;
        RECT 298.805 58.795 299.085 59.075 ;
        RECT 297.385 58.135 297.665 58.415 ;
        RECT 298.805 58.135 299.085 58.415 ;
        RECT 297.385 57.475 297.665 57.755 ;
        RECT 298.805 57.475 299.085 57.755 ;
        RECT 297.385 56.815 297.665 57.095 ;
        RECT 298.805 56.815 299.085 57.095 ;
        RECT 297.385 56.155 297.665 56.435 ;
        RECT 298.805 56.155 299.085 56.435 ;
        RECT 297.385 55.495 297.665 55.775 ;
        RECT 298.805 55.495 299.085 55.775 ;
        RECT 297.385 54.835 297.665 55.115 ;
        RECT 298.805 54.835 299.085 55.115 ;
        RECT 297.385 54.175 297.665 54.455 ;
        RECT 298.805 54.175 299.085 54.455 ;
        RECT 297.385 53.515 297.665 53.795 ;
        RECT 298.805 53.515 299.085 53.795 ;
        RECT 297.385 52.855 297.665 53.135 ;
        RECT 298.805 52.855 299.085 53.135 ;
        RECT 297.385 52.195 297.665 52.475 ;
        RECT 298.805 52.195 299.085 52.475 ;
        RECT 297.385 51.535 297.665 51.815 ;
        RECT 298.805 51.535 299.085 51.815 ;
        RECT 297.385 50.875 297.665 51.155 ;
        RECT 298.805 50.875 299.085 51.155 ;
        RECT 297.385 50.215 297.665 50.495 ;
        RECT 298.805 50.215 299.085 50.495 ;
        RECT 303.290 47.855 303.570 48.135 ;
        RECT 303.950 47.855 304.230 48.135 ;
        RECT 304.610 47.855 304.890 48.135 ;
        RECT 303.290 47.195 303.570 47.475 ;
        RECT 303.950 47.195 304.230 47.475 ;
        RECT 304.610 47.195 304.890 47.475 ;
        RECT 303.290 46.535 303.570 46.815 ;
        RECT 303.950 46.535 304.230 46.815 ;
        RECT 304.610 46.535 304.890 46.815 ;
        RECT 291.595 39.755 291.875 40.035 ;
        RECT 292.255 39.755 292.535 40.035 ;
        RECT 292.915 39.755 293.195 40.035 ;
        RECT 291.595 39.095 291.875 39.375 ;
        RECT 292.255 39.095 292.535 39.375 ;
        RECT 292.915 39.095 293.195 39.375 ;
        RECT 291.595 38.435 291.875 38.715 ;
        RECT 292.255 38.435 292.535 38.715 ;
        RECT 292.915 38.435 293.195 38.715 ;
        RECT 291.595 30.355 291.875 30.635 ;
        RECT 292.255 30.355 292.535 30.635 ;
        RECT 292.915 30.355 293.195 30.635 ;
        RECT 291.595 29.695 291.875 29.975 ;
        RECT 292.255 29.695 292.535 29.975 ;
        RECT 292.915 29.695 293.195 29.975 ;
        RECT 291.595 29.035 291.875 29.315 ;
        RECT 292.255 29.035 292.535 29.315 ;
        RECT 292.915 29.035 293.195 29.315 ;
        RECT 303.290 22.255 303.570 22.535 ;
        RECT 303.950 22.255 304.230 22.535 ;
        RECT 304.610 22.255 304.890 22.535 ;
        RECT 303.290 21.595 303.570 21.875 ;
        RECT 303.950 21.595 304.230 21.875 ;
        RECT 304.610 21.595 304.890 21.875 ;
        RECT 303.290 20.935 303.570 21.215 ;
        RECT 303.950 20.935 304.230 21.215 ;
        RECT 304.610 20.935 304.890 21.215 ;
        RECT 229.200 4.740 229.480 5.020 ;
        RECT 229.860 4.740 230.140 5.020 ;
        RECT 230.520 4.740 230.800 5.020 ;
        RECT 231.440 4.740 231.720 5.020 ;
        RECT 232.100 4.740 232.380 5.020 ;
        RECT 232.760 4.740 233.040 5.020 ;
        RECT 233.680 4.740 233.960 5.020 ;
        RECT 234.340 4.740 234.620 5.020 ;
        RECT 235.000 4.740 235.280 5.020 ;
        RECT 235.920 4.740 236.200 5.020 ;
        RECT 236.580 4.740 236.860 5.020 ;
        RECT 237.240 4.740 237.520 5.020 ;
        RECT 238.280 4.740 238.560 5.020 ;
        RECT 239.280 4.740 239.560 5.020 ;
        RECT 239.940 4.740 240.220 5.020 ;
        RECT 240.600 4.740 240.880 5.020 ;
        RECT 241.520 4.740 241.800 5.020 ;
        RECT 242.180 4.740 242.460 5.020 ;
        RECT 242.840 4.740 243.120 5.020 ;
        RECT 243.760 4.740 244.040 5.020 ;
        RECT 244.420 4.740 244.700 5.020 ;
        RECT 245.080 4.740 245.360 5.020 ;
        RECT 246.000 4.740 246.280 5.020 ;
        RECT 246.660 4.740 246.940 5.020 ;
        RECT 247.320 4.740 247.600 5.020 ;
        RECT 248.240 4.740 248.520 5.020 ;
        RECT 248.900 4.740 249.180 5.020 ;
        RECT 249.560 4.740 249.840 5.020 ;
        RECT 250.480 4.740 250.760 5.020 ;
        RECT 251.140 4.740 251.420 5.020 ;
        RECT 251.800 4.740 252.080 5.020 ;
        RECT 252.720 4.740 253.000 5.020 ;
        RECT 253.380 4.740 253.660 5.020 ;
        RECT 254.040 4.740 254.320 5.020 ;
        RECT 254.960 4.740 255.240 5.020 ;
        RECT 255.620 4.740 255.900 5.020 ;
        RECT 256.280 4.740 256.560 5.020 ;
        RECT 257.200 4.740 257.480 5.020 ;
        RECT 257.860 4.740 258.140 5.020 ;
        RECT 258.520 4.740 258.800 5.020 ;
        RECT 259.560 4.740 259.840 5.020 ;
        RECT 260.560 4.740 260.840 5.020 ;
        RECT 261.220 4.740 261.500 5.020 ;
        RECT 261.880 4.740 262.160 5.020 ;
        RECT 262.800 4.740 263.080 5.020 ;
        RECT 263.460 4.740 263.740 5.020 ;
        RECT 264.120 4.740 264.400 5.020 ;
        RECT 265.040 4.740 265.320 5.020 ;
        RECT 265.700 4.740 265.980 5.020 ;
        RECT 266.360 4.740 266.640 5.020 ;
        RECT 267.380 4.740 267.660 5.020 ;
        RECT 268.040 4.740 268.320 5.020 ;
        RECT 268.700 4.740 268.980 5.020 ;
        RECT 309.095 58.795 309.375 59.075 ;
        RECT 309.095 58.135 309.375 58.415 ;
        RECT 309.095 57.475 309.375 57.755 ;
        RECT 309.095 56.815 309.375 57.095 ;
        RECT 309.095 56.155 309.375 56.435 ;
        RECT 309.095 55.495 309.375 55.775 ;
        RECT 309.095 54.835 309.375 55.115 ;
        RECT 309.095 54.175 309.375 54.455 ;
        RECT 309.095 53.515 309.375 53.795 ;
        RECT 309.095 52.855 309.375 53.135 ;
        RECT 309.095 52.195 309.375 52.475 ;
        RECT 309.095 51.535 309.375 51.815 ;
        RECT 309.095 50.875 309.375 51.155 ;
        RECT 309.095 50.215 309.375 50.495 ;
        RECT 319.380 58.795 319.660 59.075 ;
        RECT 319.380 58.135 319.660 58.415 ;
        RECT 319.380 57.475 319.660 57.755 ;
        RECT 319.380 56.815 319.660 57.095 ;
        RECT 319.380 56.155 319.660 56.435 ;
        RECT 319.380 55.495 319.660 55.775 ;
        RECT 319.380 54.835 319.660 55.115 ;
        RECT 319.380 54.175 319.660 54.455 ;
        RECT 319.380 53.515 319.660 53.795 ;
        RECT 319.380 52.855 319.660 53.135 ;
        RECT 319.380 52.195 319.660 52.475 ;
        RECT 319.380 51.535 319.660 51.815 ;
        RECT 319.380 50.875 319.660 51.155 ;
        RECT 319.380 50.215 319.660 50.495 ;
        RECT 313.590 45.155 313.870 45.435 ;
        RECT 314.250 45.155 314.530 45.435 ;
        RECT 314.910 45.155 315.190 45.435 ;
        RECT 313.590 44.495 313.870 44.775 ;
        RECT 314.250 44.495 314.530 44.775 ;
        RECT 314.910 44.495 315.190 44.775 ;
        RECT 313.590 43.835 313.870 44.115 ;
        RECT 314.250 43.835 314.530 44.115 ;
        RECT 314.910 43.835 315.190 44.115 ;
        RECT 323.865 42.455 324.145 42.735 ;
        RECT 324.525 42.455 324.805 42.735 ;
        RECT 325.185 42.455 325.465 42.735 ;
        RECT 323.865 41.795 324.145 42.075 ;
        RECT 324.525 41.795 324.805 42.075 ;
        RECT 325.185 41.795 325.465 42.075 ;
        RECT 323.865 41.135 324.145 41.415 ;
        RECT 324.525 41.135 324.805 41.415 ;
        RECT 325.185 41.135 325.465 41.415 ;
        RECT 323.865 27.655 324.145 27.935 ;
        RECT 324.525 27.655 324.805 27.935 ;
        RECT 325.185 27.655 325.465 27.935 ;
        RECT 323.865 26.995 324.145 27.275 ;
        RECT 324.525 26.995 324.805 27.275 ;
        RECT 325.185 26.995 325.465 27.275 ;
        RECT 323.865 26.335 324.145 26.615 ;
        RECT 324.525 26.335 324.805 26.615 ;
        RECT 325.185 26.335 325.465 26.615 ;
        RECT 313.590 24.955 313.870 25.235 ;
        RECT 314.250 24.955 314.530 25.235 ;
        RECT 314.910 24.955 315.190 25.235 ;
        RECT 313.590 24.295 313.870 24.575 ;
        RECT 314.250 24.295 314.530 24.575 ;
        RECT 314.910 24.295 315.190 24.575 ;
        RECT 313.590 23.635 313.870 23.915 ;
        RECT 314.250 23.635 314.530 23.915 ;
        RECT 314.910 23.635 315.190 23.915 ;
        RECT 329.670 58.795 329.950 59.075 ;
        RECT 329.670 58.135 329.950 58.415 ;
        RECT 329.670 57.475 329.950 57.755 ;
        RECT 329.670 56.815 329.950 57.095 ;
        RECT 329.670 56.155 329.950 56.435 ;
        RECT 329.670 55.495 329.950 55.775 ;
        RECT 329.670 54.835 329.950 55.115 ;
        RECT 329.670 54.175 329.950 54.455 ;
        RECT 329.670 53.515 329.950 53.795 ;
        RECT 329.670 52.855 329.950 53.135 ;
        RECT 329.670 52.195 329.950 52.475 ;
        RECT 329.670 51.535 329.950 51.815 ;
        RECT 329.670 50.875 329.950 51.155 ;
        RECT 329.670 50.215 329.950 50.495 ;
        RECT 339.955 58.795 340.235 59.075 ;
        RECT 341.375 58.795 341.655 59.075 ;
        RECT 339.955 58.135 340.235 58.415 ;
        RECT 341.375 58.135 341.655 58.415 ;
        RECT 339.955 57.475 340.235 57.755 ;
        RECT 341.375 57.475 341.655 57.755 ;
        RECT 339.955 56.815 340.235 57.095 ;
        RECT 341.375 56.815 341.655 57.095 ;
        RECT 339.955 56.155 340.235 56.435 ;
        RECT 341.375 56.155 341.655 56.435 ;
        RECT 339.955 55.495 340.235 55.775 ;
        RECT 341.375 55.495 341.655 55.775 ;
        RECT 339.955 54.835 340.235 55.115 ;
        RECT 341.375 54.835 341.655 55.115 ;
        RECT 339.955 54.175 340.235 54.455 ;
        RECT 341.375 54.175 341.655 54.455 ;
        RECT 339.955 53.515 340.235 53.795 ;
        RECT 341.375 53.515 341.655 53.795 ;
        RECT 339.955 52.855 340.235 53.135 ;
        RECT 341.375 52.855 341.655 53.135 ;
        RECT 339.955 52.195 340.235 52.475 ;
        RECT 341.375 52.195 341.655 52.475 ;
        RECT 339.955 51.535 340.235 51.815 ;
        RECT 341.375 51.535 341.655 51.815 ;
        RECT 339.955 50.875 340.235 51.155 ;
        RECT 341.375 50.875 341.655 51.155 ;
        RECT 339.955 50.215 340.235 50.495 ;
        RECT 341.375 50.215 341.655 50.495 ;
        RECT 345.860 47.855 346.140 48.135 ;
        RECT 346.520 47.855 346.800 48.135 ;
        RECT 347.180 47.855 347.460 48.135 ;
        RECT 345.860 47.195 346.140 47.475 ;
        RECT 346.520 47.195 346.800 47.475 ;
        RECT 347.180 47.195 347.460 47.475 ;
        RECT 345.860 46.535 346.140 46.815 ;
        RECT 346.520 46.535 346.800 46.815 ;
        RECT 347.180 46.535 347.460 46.815 ;
        RECT 334.165 39.755 334.445 40.035 ;
        RECT 334.825 39.755 335.105 40.035 ;
        RECT 335.485 39.755 335.765 40.035 ;
        RECT 334.165 39.095 334.445 39.375 ;
        RECT 334.825 39.095 335.105 39.375 ;
        RECT 335.485 39.095 335.765 39.375 ;
        RECT 334.165 38.435 334.445 38.715 ;
        RECT 334.825 38.435 335.105 38.715 ;
        RECT 335.485 38.435 335.765 38.715 ;
        RECT 334.165 30.355 334.445 30.635 ;
        RECT 334.825 30.355 335.105 30.635 ;
        RECT 335.485 30.355 335.765 30.635 ;
        RECT 334.165 29.695 334.445 29.975 ;
        RECT 334.825 29.695 335.105 29.975 ;
        RECT 335.485 29.695 335.765 29.975 ;
        RECT 334.165 29.035 334.445 29.315 ;
        RECT 334.825 29.035 335.105 29.315 ;
        RECT 335.485 29.035 335.765 29.315 ;
        RECT 345.860 22.255 346.140 22.535 ;
        RECT 346.520 22.255 346.800 22.535 ;
        RECT 347.180 22.255 347.460 22.535 ;
        RECT 345.860 21.595 346.140 21.875 ;
        RECT 346.520 21.595 346.800 21.875 ;
        RECT 347.180 21.595 347.460 21.875 ;
        RECT 345.860 20.935 346.140 21.215 ;
        RECT 346.520 20.935 346.800 21.215 ;
        RECT 347.180 20.935 347.460 21.215 ;
        RECT 270.640 4.740 270.920 5.020 ;
        RECT 271.300 4.740 271.580 5.020 ;
        RECT 271.960 4.740 272.240 5.020 ;
        RECT 272.880 4.740 273.160 5.020 ;
        RECT 273.540 4.740 273.820 5.020 ;
        RECT 274.200 4.740 274.480 5.020 ;
        RECT 275.120 4.740 275.400 5.020 ;
        RECT 275.780 4.740 276.060 5.020 ;
        RECT 276.440 4.740 276.720 5.020 ;
        RECT 277.360 4.740 277.640 5.020 ;
        RECT 278.020 4.740 278.300 5.020 ;
        RECT 278.680 4.740 278.960 5.020 ;
        RECT 279.720 4.740 280.000 5.020 ;
        RECT 280.720 4.740 281.000 5.020 ;
        RECT 281.380 4.740 281.660 5.020 ;
        RECT 282.040 4.740 282.320 5.020 ;
        RECT 282.960 4.740 283.240 5.020 ;
        RECT 283.620 4.740 283.900 5.020 ;
        RECT 284.280 4.740 284.560 5.020 ;
        RECT 285.200 4.740 285.480 5.020 ;
        RECT 285.860 4.740 286.140 5.020 ;
        RECT 286.520 4.740 286.800 5.020 ;
        RECT 287.440 4.740 287.720 5.020 ;
        RECT 288.100 4.740 288.380 5.020 ;
        RECT 288.760 4.740 289.040 5.020 ;
        RECT 289.680 4.740 289.960 5.020 ;
        RECT 290.340 4.740 290.620 5.020 ;
        RECT 291.000 4.740 291.280 5.020 ;
        RECT 291.920 4.740 292.200 5.020 ;
        RECT 292.580 4.740 292.860 5.020 ;
        RECT 293.240 4.740 293.520 5.020 ;
        RECT 294.160 4.740 294.440 5.020 ;
        RECT 294.820 4.740 295.100 5.020 ;
        RECT 295.480 4.740 295.760 5.020 ;
        RECT 296.400 4.740 296.680 5.020 ;
        RECT 297.060 4.740 297.340 5.020 ;
        RECT 297.720 4.740 298.000 5.020 ;
        RECT 298.640 4.740 298.920 5.020 ;
        RECT 299.300 4.740 299.580 5.020 ;
        RECT 299.960 4.740 300.240 5.020 ;
        RECT 301.000 4.740 301.280 5.020 ;
        RECT 302.000 4.740 302.280 5.020 ;
        RECT 302.660 4.740 302.940 5.020 ;
        RECT 303.320 4.740 303.600 5.020 ;
        RECT 304.240 4.740 304.520 5.020 ;
        RECT 304.900 4.740 305.180 5.020 ;
        RECT 305.560 4.740 305.840 5.020 ;
        RECT 306.480 4.740 306.760 5.020 ;
        RECT 307.140 4.740 307.420 5.020 ;
        RECT 307.800 4.740 308.080 5.020 ;
        RECT 308.720 4.740 309.000 5.020 ;
        RECT 309.380 4.740 309.660 5.020 ;
        RECT 310.040 4.740 310.320 5.020 ;
        RECT 311.060 4.740 311.340 5.020 ;
        RECT 311.720 4.740 312.000 5.020 ;
        RECT 312.380 4.740 312.660 5.020 ;
        RECT 351.665 58.795 351.945 59.075 ;
        RECT 351.665 58.135 351.945 58.415 ;
        RECT 351.665 57.475 351.945 57.755 ;
        RECT 351.665 56.815 351.945 57.095 ;
        RECT 351.665 56.155 351.945 56.435 ;
        RECT 351.665 55.495 351.945 55.775 ;
        RECT 351.665 54.835 351.945 55.115 ;
        RECT 351.665 54.175 351.945 54.455 ;
        RECT 351.665 53.515 351.945 53.795 ;
        RECT 351.665 52.855 351.945 53.135 ;
        RECT 351.665 52.195 351.945 52.475 ;
        RECT 351.665 51.535 351.945 51.815 ;
        RECT 351.665 50.875 351.945 51.155 ;
        RECT 351.665 50.215 351.945 50.495 ;
        RECT 361.950 58.795 362.230 59.075 ;
        RECT 361.950 58.135 362.230 58.415 ;
        RECT 361.950 57.475 362.230 57.755 ;
        RECT 361.950 56.815 362.230 57.095 ;
        RECT 361.950 56.155 362.230 56.435 ;
        RECT 361.950 55.495 362.230 55.775 ;
        RECT 361.950 54.835 362.230 55.115 ;
        RECT 361.950 54.175 362.230 54.455 ;
        RECT 361.950 53.515 362.230 53.795 ;
        RECT 361.950 52.855 362.230 53.135 ;
        RECT 361.950 52.195 362.230 52.475 ;
        RECT 361.950 51.535 362.230 51.815 ;
        RECT 361.950 50.875 362.230 51.155 ;
        RECT 361.950 50.215 362.230 50.495 ;
        RECT 356.160 45.155 356.440 45.435 ;
        RECT 356.820 45.155 357.100 45.435 ;
        RECT 357.480 45.155 357.760 45.435 ;
        RECT 356.160 44.495 356.440 44.775 ;
        RECT 356.820 44.495 357.100 44.775 ;
        RECT 357.480 44.495 357.760 44.775 ;
        RECT 356.160 43.835 356.440 44.115 ;
        RECT 356.820 43.835 357.100 44.115 ;
        RECT 357.480 43.835 357.760 44.115 ;
        RECT 366.435 42.455 366.715 42.735 ;
        RECT 367.095 42.455 367.375 42.735 ;
        RECT 367.755 42.455 368.035 42.735 ;
        RECT 366.435 41.795 366.715 42.075 ;
        RECT 367.095 41.795 367.375 42.075 ;
        RECT 367.755 41.795 368.035 42.075 ;
        RECT 366.435 41.135 366.715 41.415 ;
        RECT 367.095 41.135 367.375 41.415 ;
        RECT 367.755 41.135 368.035 41.415 ;
        RECT 366.435 27.655 366.715 27.935 ;
        RECT 367.095 27.655 367.375 27.935 ;
        RECT 367.755 27.655 368.035 27.935 ;
        RECT 366.435 26.995 366.715 27.275 ;
        RECT 367.095 26.995 367.375 27.275 ;
        RECT 367.755 26.995 368.035 27.275 ;
        RECT 366.435 26.335 366.715 26.615 ;
        RECT 367.095 26.335 367.375 26.615 ;
        RECT 367.755 26.335 368.035 26.615 ;
        RECT 356.160 24.955 356.440 25.235 ;
        RECT 356.820 24.955 357.100 25.235 ;
        RECT 357.480 24.955 357.760 25.235 ;
        RECT 356.160 24.295 356.440 24.575 ;
        RECT 356.820 24.295 357.100 24.575 ;
        RECT 357.480 24.295 357.760 24.575 ;
        RECT 356.160 23.635 356.440 23.915 ;
        RECT 356.820 23.635 357.100 23.915 ;
        RECT 357.480 23.635 357.760 23.915 ;
        RECT 372.240 58.795 372.520 59.075 ;
        RECT 372.240 58.135 372.520 58.415 ;
        RECT 372.240 57.475 372.520 57.755 ;
        RECT 372.240 56.815 372.520 57.095 ;
        RECT 372.240 56.155 372.520 56.435 ;
        RECT 372.240 55.495 372.520 55.775 ;
        RECT 372.240 54.835 372.520 55.115 ;
        RECT 372.240 54.175 372.520 54.455 ;
        RECT 372.240 53.515 372.520 53.795 ;
        RECT 372.240 52.855 372.520 53.135 ;
        RECT 372.240 52.195 372.520 52.475 ;
        RECT 372.240 51.535 372.520 51.815 ;
        RECT 372.240 50.875 372.520 51.155 ;
        RECT 372.240 50.215 372.520 50.495 ;
        RECT 382.525 58.795 382.805 59.075 ;
        RECT 383.945 58.795 384.225 59.075 ;
        RECT 382.525 58.135 382.805 58.415 ;
        RECT 383.945 58.135 384.225 58.415 ;
        RECT 382.525 57.475 382.805 57.755 ;
        RECT 383.945 57.475 384.225 57.755 ;
        RECT 382.525 56.815 382.805 57.095 ;
        RECT 383.945 56.815 384.225 57.095 ;
        RECT 382.525 56.155 382.805 56.435 ;
        RECT 383.945 56.155 384.225 56.435 ;
        RECT 382.525 55.495 382.805 55.775 ;
        RECT 383.945 55.495 384.225 55.775 ;
        RECT 382.525 54.835 382.805 55.115 ;
        RECT 383.945 54.835 384.225 55.115 ;
        RECT 382.525 54.175 382.805 54.455 ;
        RECT 383.945 54.175 384.225 54.455 ;
        RECT 382.525 53.515 382.805 53.795 ;
        RECT 383.945 53.515 384.225 53.795 ;
        RECT 382.525 52.855 382.805 53.135 ;
        RECT 383.945 52.855 384.225 53.135 ;
        RECT 382.525 52.195 382.805 52.475 ;
        RECT 383.945 52.195 384.225 52.475 ;
        RECT 382.525 51.535 382.805 51.815 ;
        RECT 383.945 51.535 384.225 51.815 ;
        RECT 382.525 50.875 382.805 51.155 ;
        RECT 383.945 50.875 384.225 51.155 ;
        RECT 382.525 50.215 382.805 50.495 ;
        RECT 383.945 50.215 384.225 50.495 ;
        RECT 388.430 47.855 388.710 48.135 ;
        RECT 389.090 47.855 389.370 48.135 ;
        RECT 389.750 47.855 390.030 48.135 ;
        RECT 388.430 47.195 388.710 47.475 ;
        RECT 389.090 47.195 389.370 47.475 ;
        RECT 389.750 47.195 390.030 47.475 ;
        RECT 388.430 46.535 388.710 46.815 ;
        RECT 389.090 46.535 389.370 46.815 ;
        RECT 389.750 46.535 390.030 46.815 ;
        RECT 376.735 39.755 377.015 40.035 ;
        RECT 377.395 39.755 377.675 40.035 ;
        RECT 378.055 39.755 378.335 40.035 ;
        RECT 376.735 39.095 377.015 39.375 ;
        RECT 377.395 39.095 377.675 39.375 ;
        RECT 378.055 39.095 378.335 39.375 ;
        RECT 376.735 38.435 377.015 38.715 ;
        RECT 377.395 38.435 377.675 38.715 ;
        RECT 378.055 38.435 378.335 38.715 ;
        RECT 376.735 30.355 377.015 30.635 ;
        RECT 377.395 30.355 377.675 30.635 ;
        RECT 378.055 30.355 378.335 30.635 ;
        RECT 376.735 29.695 377.015 29.975 ;
        RECT 377.395 29.695 377.675 29.975 ;
        RECT 378.055 29.695 378.335 29.975 ;
        RECT 376.735 29.035 377.015 29.315 ;
        RECT 377.395 29.035 377.675 29.315 ;
        RECT 378.055 29.035 378.335 29.315 ;
        RECT 388.430 22.255 388.710 22.535 ;
        RECT 389.090 22.255 389.370 22.535 ;
        RECT 389.750 22.255 390.030 22.535 ;
        RECT 388.430 21.595 388.710 21.875 ;
        RECT 389.090 21.595 389.370 21.875 ;
        RECT 389.750 21.595 390.030 21.875 ;
        RECT 388.430 20.935 388.710 21.215 ;
        RECT 389.090 20.935 389.370 21.215 ;
        RECT 389.750 20.935 390.030 21.215 ;
        RECT 314.320 4.740 314.600 5.020 ;
        RECT 314.980 4.740 315.260 5.020 ;
        RECT 315.640 4.740 315.920 5.020 ;
        RECT 316.560 4.740 316.840 5.020 ;
        RECT 317.220 4.740 317.500 5.020 ;
        RECT 317.880 4.740 318.160 5.020 ;
        RECT 318.800 4.740 319.080 5.020 ;
        RECT 319.460 4.740 319.740 5.020 ;
        RECT 320.120 4.740 320.400 5.020 ;
        RECT 321.160 4.740 321.440 5.020 ;
        RECT 322.160 4.740 322.440 5.020 ;
        RECT 322.820 4.740 323.100 5.020 ;
        RECT 323.480 4.740 323.760 5.020 ;
        RECT 324.400 4.740 324.680 5.020 ;
        RECT 325.060 4.740 325.340 5.020 ;
        RECT 325.720 4.740 326.000 5.020 ;
        RECT 326.640 4.740 326.920 5.020 ;
        RECT 327.300 4.740 327.580 5.020 ;
        RECT 327.960 4.740 328.240 5.020 ;
        RECT 328.880 4.740 329.160 5.020 ;
        RECT 329.540 4.740 329.820 5.020 ;
        RECT 330.200 4.740 330.480 5.020 ;
        RECT 331.120 4.740 331.400 5.020 ;
        RECT 331.780 4.740 332.060 5.020 ;
        RECT 332.440 4.740 332.720 5.020 ;
        RECT 333.360 4.740 333.640 5.020 ;
        RECT 334.020 4.740 334.300 5.020 ;
        RECT 334.680 4.740 334.960 5.020 ;
        RECT 335.600 4.740 335.880 5.020 ;
        RECT 336.260 4.740 336.540 5.020 ;
        RECT 336.920 4.740 337.200 5.020 ;
        RECT 337.840 4.740 338.120 5.020 ;
        RECT 338.500 4.740 338.780 5.020 ;
        RECT 339.160 4.740 339.440 5.020 ;
        RECT 340.080 4.740 340.360 5.020 ;
        RECT 340.740 4.740 341.020 5.020 ;
        RECT 341.400 4.740 341.680 5.020 ;
        RECT 342.440 4.740 342.720 5.020 ;
        RECT 343.440 4.740 343.720 5.020 ;
        RECT 344.100 4.740 344.380 5.020 ;
        RECT 344.760 4.740 345.040 5.020 ;
        RECT 345.680 4.740 345.960 5.020 ;
        RECT 346.340 4.740 346.620 5.020 ;
        RECT 347.000 4.740 347.280 5.020 ;
        RECT 347.920 4.740 348.200 5.020 ;
        RECT 348.580 4.740 348.860 5.020 ;
        RECT 349.240 4.740 349.520 5.020 ;
        RECT 350.160 4.740 350.440 5.020 ;
        RECT 350.820 4.740 351.100 5.020 ;
        RECT 351.480 4.740 351.760 5.020 ;
        RECT 352.500 4.740 352.780 5.020 ;
        RECT 353.160 4.740 353.440 5.020 ;
        RECT 353.820 4.740 354.100 5.020 ;
        RECT 394.235 58.795 394.515 59.075 ;
        RECT 394.235 58.135 394.515 58.415 ;
        RECT 394.235 57.475 394.515 57.755 ;
        RECT 394.235 56.815 394.515 57.095 ;
        RECT 394.235 56.155 394.515 56.435 ;
        RECT 394.235 55.495 394.515 55.775 ;
        RECT 394.235 54.835 394.515 55.115 ;
        RECT 394.235 54.175 394.515 54.455 ;
        RECT 394.235 53.515 394.515 53.795 ;
        RECT 394.235 52.855 394.515 53.135 ;
        RECT 394.235 52.195 394.515 52.475 ;
        RECT 394.235 51.535 394.515 51.815 ;
        RECT 394.235 50.875 394.515 51.155 ;
        RECT 394.235 50.215 394.515 50.495 ;
        RECT 404.520 58.795 404.800 59.075 ;
        RECT 404.520 58.135 404.800 58.415 ;
        RECT 404.520 57.475 404.800 57.755 ;
        RECT 404.520 56.815 404.800 57.095 ;
        RECT 404.520 56.155 404.800 56.435 ;
        RECT 404.520 55.495 404.800 55.775 ;
        RECT 404.520 54.835 404.800 55.115 ;
        RECT 404.520 54.175 404.800 54.455 ;
        RECT 404.520 53.515 404.800 53.795 ;
        RECT 404.520 52.855 404.800 53.135 ;
        RECT 404.520 52.195 404.800 52.475 ;
        RECT 404.520 51.535 404.800 51.815 ;
        RECT 404.520 50.875 404.800 51.155 ;
        RECT 404.520 50.215 404.800 50.495 ;
        RECT 398.730 45.155 399.010 45.435 ;
        RECT 399.390 45.155 399.670 45.435 ;
        RECT 400.050 45.155 400.330 45.435 ;
        RECT 398.730 44.495 399.010 44.775 ;
        RECT 399.390 44.495 399.670 44.775 ;
        RECT 400.050 44.495 400.330 44.775 ;
        RECT 398.730 43.835 399.010 44.115 ;
        RECT 399.390 43.835 399.670 44.115 ;
        RECT 400.050 43.835 400.330 44.115 ;
        RECT 409.005 42.455 409.285 42.735 ;
        RECT 409.665 42.455 409.945 42.735 ;
        RECT 410.325 42.455 410.605 42.735 ;
        RECT 409.005 41.795 409.285 42.075 ;
        RECT 409.665 41.795 409.945 42.075 ;
        RECT 410.325 41.795 410.605 42.075 ;
        RECT 409.005 41.135 409.285 41.415 ;
        RECT 409.665 41.135 409.945 41.415 ;
        RECT 410.325 41.135 410.605 41.415 ;
        RECT 409.005 27.655 409.285 27.935 ;
        RECT 409.665 27.655 409.945 27.935 ;
        RECT 410.325 27.655 410.605 27.935 ;
        RECT 409.005 26.995 409.285 27.275 ;
        RECT 409.665 26.995 409.945 27.275 ;
        RECT 410.325 26.995 410.605 27.275 ;
        RECT 409.005 26.335 409.285 26.615 ;
        RECT 409.665 26.335 409.945 26.615 ;
        RECT 410.325 26.335 410.605 26.615 ;
        RECT 398.730 24.955 399.010 25.235 ;
        RECT 399.390 24.955 399.670 25.235 ;
        RECT 400.050 24.955 400.330 25.235 ;
        RECT 398.730 24.295 399.010 24.575 ;
        RECT 399.390 24.295 399.670 24.575 ;
        RECT 400.050 24.295 400.330 24.575 ;
        RECT 398.730 23.635 399.010 23.915 ;
        RECT 399.390 23.635 399.670 23.915 ;
        RECT 400.050 23.635 400.330 23.915 ;
        RECT 414.810 58.795 415.090 59.075 ;
        RECT 414.810 58.135 415.090 58.415 ;
        RECT 414.810 57.475 415.090 57.755 ;
        RECT 414.810 56.815 415.090 57.095 ;
        RECT 414.810 56.155 415.090 56.435 ;
        RECT 414.810 55.495 415.090 55.775 ;
        RECT 414.810 54.835 415.090 55.115 ;
        RECT 414.810 54.175 415.090 54.455 ;
        RECT 414.810 53.515 415.090 53.795 ;
        RECT 414.810 52.855 415.090 53.135 ;
        RECT 414.810 52.195 415.090 52.475 ;
        RECT 414.810 51.535 415.090 51.815 ;
        RECT 414.810 50.875 415.090 51.155 ;
        RECT 414.810 50.215 415.090 50.495 ;
        RECT 425.095 58.795 425.375 59.075 ;
        RECT 426.515 58.795 426.795 59.075 ;
        RECT 425.095 58.135 425.375 58.415 ;
        RECT 426.515 58.135 426.795 58.415 ;
        RECT 425.095 57.475 425.375 57.755 ;
        RECT 426.515 57.475 426.795 57.755 ;
        RECT 425.095 56.815 425.375 57.095 ;
        RECT 426.515 56.815 426.795 57.095 ;
        RECT 425.095 56.155 425.375 56.435 ;
        RECT 426.515 56.155 426.795 56.435 ;
        RECT 425.095 55.495 425.375 55.775 ;
        RECT 426.515 55.495 426.795 55.775 ;
        RECT 425.095 54.835 425.375 55.115 ;
        RECT 426.515 54.835 426.795 55.115 ;
        RECT 425.095 54.175 425.375 54.455 ;
        RECT 426.515 54.175 426.795 54.455 ;
        RECT 425.095 53.515 425.375 53.795 ;
        RECT 426.515 53.515 426.795 53.795 ;
        RECT 425.095 52.855 425.375 53.135 ;
        RECT 426.515 52.855 426.795 53.135 ;
        RECT 425.095 52.195 425.375 52.475 ;
        RECT 426.515 52.195 426.795 52.475 ;
        RECT 425.095 51.535 425.375 51.815 ;
        RECT 426.515 51.535 426.795 51.815 ;
        RECT 425.095 50.875 425.375 51.155 ;
        RECT 426.515 50.875 426.795 51.155 ;
        RECT 425.095 50.215 425.375 50.495 ;
        RECT 426.515 50.215 426.795 50.495 ;
        RECT 431.000 47.855 431.280 48.135 ;
        RECT 431.660 47.855 431.940 48.135 ;
        RECT 432.320 47.855 432.600 48.135 ;
        RECT 431.000 47.195 431.280 47.475 ;
        RECT 431.660 47.195 431.940 47.475 ;
        RECT 432.320 47.195 432.600 47.475 ;
        RECT 431.000 46.535 431.280 46.815 ;
        RECT 431.660 46.535 431.940 46.815 ;
        RECT 432.320 46.535 432.600 46.815 ;
        RECT 419.305 39.755 419.585 40.035 ;
        RECT 419.965 39.755 420.245 40.035 ;
        RECT 420.625 39.755 420.905 40.035 ;
        RECT 419.305 39.095 419.585 39.375 ;
        RECT 419.965 39.095 420.245 39.375 ;
        RECT 420.625 39.095 420.905 39.375 ;
        RECT 419.305 38.435 419.585 38.715 ;
        RECT 419.965 38.435 420.245 38.715 ;
        RECT 420.625 38.435 420.905 38.715 ;
        RECT 419.305 30.355 419.585 30.635 ;
        RECT 419.965 30.355 420.245 30.635 ;
        RECT 420.625 30.355 420.905 30.635 ;
        RECT 419.305 29.695 419.585 29.975 ;
        RECT 419.965 29.695 420.245 29.975 ;
        RECT 420.625 29.695 420.905 29.975 ;
        RECT 419.305 29.035 419.585 29.315 ;
        RECT 419.965 29.035 420.245 29.315 ;
        RECT 420.625 29.035 420.905 29.315 ;
        RECT 431.000 22.255 431.280 22.535 ;
        RECT 431.660 22.255 431.940 22.535 ;
        RECT 432.320 22.255 432.600 22.535 ;
        RECT 431.000 21.595 431.280 21.875 ;
        RECT 431.660 21.595 431.940 21.875 ;
        RECT 432.320 21.595 432.600 21.875 ;
        RECT 431.000 20.935 431.280 21.215 ;
        RECT 431.660 20.935 431.940 21.215 ;
        RECT 432.320 20.935 432.600 21.215 ;
        RECT 355.760 4.740 356.040 5.020 ;
        RECT 356.420 4.740 356.700 5.020 ;
        RECT 357.080 4.740 357.360 5.020 ;
        RECT 358.000 4.740 358.280 5.020 ;
        RECT 358.660 4.740 358.940 5.020 ;
        RECT 359.320 4.740 359.600 5.020 ;
        RECT 360.240 4.740 360.520 5.020 ;
        RECT 360.900 4.740 361.180 5.020 ;
        RECT 361.560 4.740 361.840 5.020 ;
        RECT 362.600 4.740 362.880 5.020 ;
        RECT 363.600 4.740 363.880 5.020 ;
        RECT 364.260 4.740 364.540 5.020 ;
        RECT 364.920 4.740 365.200 5.020 ;
        RECT 365.840 4.740 366.120 5.020 ;
        RECT 366.500 4.740 366.780 5.020 ;
        RECT 367.160 4.740 367.440 5.020 ;
        RECT 368.080 4.740 368.360 5.020 ;
        RECT 368.740 4.740 369.020 5.020 ;
        RECT 369.400 4.740 369.680 5.020 ;
        RECT 370.320 4.740 370.600 5.020 ;
        RECT 370.980 4.740 371.260 5.020 ;
        RECT 371.640 4.740 371.920 5.020 ;
        RECT 372.560 4.740 372.840 5.020 ;
        RECT 373.220 4.740 373.500 5.020 ;
        RECT 373.880 4.740 374.160 5.020 ;
        RECT 374.800 4.740 375.080 5.020 ;
        RECT 375.460 4.740 375.740 5.020 ;
        RECT 376.120 4.740 376.400 5.020 ;
        RECT 377.040 4.740 377.320 5.020 ;
        RECT 377.700 4.740 377.980 5.020 ;
        RECT 378.360 4.740 378.640 5.020 ;
        RECT 379.280 4.740 379.560 5.020 ;
        RECT 379.940 4.740 380.220 5.020 ;
        RECT 380.600 4.740 380.880 5.020 ;
        RECT 381.520 4.740 381.800 5.020 ;
        RECT 382.180 4.740 382.460 5.020 ;
        RECT 382.840 4.740 383.120 5.020 ;
        RECT 383.880 4.740 384.160 5.020 ;
        RECT 384.880 4.740 385.160 5.020 ;
        RECT 385.540 4.740 385.820 5.020 ;
        RECT 386.200 4.740 386.480 5.020 ;
        RECT 387.120 4.740 387.400 5.020 ;
        RECT 387.780 4.740 388.060 5.020 ;
        RECT 388.440 4.740 388.720 5.020 ;
        RECT 389.360 4.740 389.640 5.020 ;
        RECT 390.020 4.740 390.300 5.020 ;
        RECT 390.680 4.740 390.960 5.020 ;
        RECT 391.600 4.740 391.880 5.020 ;
        RECT 392.260 4.740 392.540 5.020 ;
        RECT 392.920 4.740 393.200 5.020 ;
        RECT 393.840 4.740 394.120 5.020 ;
        RECT 394.500 4.740 394.780 5.020 ;
        RECT 395.160 4.740 395.440 5.020 ;
        RECT 396.180 4.740 396.460 5.020 ;
        RECT 396.840 4.740 397.120 5.020 ;
        RECT 397.500 4.740 397.780 5.020 ;
        RECT 436.805 58.795 437.085 59.075 ;
        RECT 436.805 58.135 437.085 58.415 ;
        RECT 436.805 57.475 437.085 57.755 ;
        RECT 436.805 56.815 437.085 57.095 ;
        RECT 436.805 56.155 437.085 56.435 ;
        RECT 436.805 55.495 437.085 55.775 ;
        RECT 436.805 54.835 437.085 55.115 ;
        RECT 436.805 54.175 437.085 54.455 ;
        RECT 436.805 53.515 437.085 53.795 ;
        RECT 436.805 52.855 437.085 53.135 ;
        RECT 436.805 52.195 437.085 52.475 ;
        RECT 436.805 51.535 437.085 51.815 ;
        RECT 436.805 50.875 437.085 51.155 ;
        RECT 436.805 50.215 437.085 50.495 ;
        RECT 447.090 58.795 447.370 59.075 ;
        RECT 447.090 58.135 447.370 58.415 ;
        RECT 447.090 57.475 447.370 57.755 ;
        RECT 447.090 56.815 447.370 57.095 ;
        RECT 447.090 56.155 447.370 56.435 ;
        RECT 447.090 55.495 447.370 55.775 ;
        RECT 447.090 54.835 447.370 55.115 ;
        RECT 447.090 54.175 447.370 54.455 ;
        RECT 447.090 53.515 447.370 53.795 ;
        RECT 447.090 52.855 447.370 53.135 ;
        RECT 447.090 52.195 447.370 52.475 ;
        RECT 447.090 51.535 447.370 51.815 ;
        RECT 447.090 50.875 447.370 51.155 ;
        RECT 447.090 50.215 447.370 50.495 ;
        RECT 441.300 45.155 441.580 45.435 ;
        RECT 441.960 45.155 442.240 45.435 ;
        RECT 442.620 45.155 442.900 45.435 ;
        RECT 441.300 44.495 441.580 44.775 ;
        RECT 441.960 44.495 442.240 44.775 ;
        RECT 442.620 44.495 442.900 44.775 ;
        RECT 441.300 43.835 441.580 44.115 ;
        RECT 441.960 43.835 442.240 44.115 ;
        RECT 442.620 43.835 442.900 44.115 ;
        RECT 451.575 42.455 451.855 42.735 ;
        RECT 452.235 42.455 452.515 42.735 ;
        RECT 452.895 42.455 453.175 42.735 ;
        RECT 451.575 41.795 451.855 42.075 ;
        RECT 452.235 41.795 452.515 42.075 ;
        RECT 452.895 41.795 453.175 42.075 ;
        RECT 451.575 41.135 451.855 41.415 ;
        RECT 452.235 41.135 452.515 41.415 ;
        RECT 452.895 41.135 453.175 41.415 ;
        RECT 451.575 27.655 451.855 27.935 ;
        RECT 452.235 27.655 452.515 27.935 ;
        RECT 452.895 27.655 453.175 27.935 ;
        RECT 451.575 26.995 451.855 27.275 ;
        RECT 452.235 26.995 452.515 27.275 ;
        RECT 452.895 26.995 453.175 27.275 ;
        RECT 451.575 26.335 451.855 26.615 ;
        RECT 452.235 26.335 452.515 26.615 ;
        RECT 452.895 26.335 453.175 26.615 ;
        RECT 441.300 24.955 441.580 25.235 ;
        RECT 441.960 24.955 442.240 25.235 ;
        RECT 442.620 24.955 442.900 25.235 ;
        RECT 441.300 24.295 441.580 24.575 ;
        RECT 441.960 24.295 442.240 24.575 ;
        RECT 442.620 24.295 442.900 24.575 ;
        RECT 441.300 23.635 441.580 23.915 ;
        RECT 441.960 23.635 442.240 23.915 ;
        RECT 442.620 23.635 442.900 23.915 ;
        RECT 457.380 58.795 457.660 59.075 ;
        RECT 457.380 58.135 457.660 58.415 ;
        RECT 457.380 57.475 457.660 57.755 ;
        RECT 457.380 56.815 457.660 57.095 ;
        RECT 457.380 56.155 457.660 56.435 ;
        RECT 457.380 55.495 457.660 55.775 ;
        RECT 457.380 54.835 457.660 55.115 ;
        RECT 457.380 54.175 457.660 54.455 ;
        RECT 457.380 53.515 457.660 53.795 ;
        RECT 457.380 52.855 457.660 53.135 ;
        RECT 457.380 52.195 457.660 52.475 ;
        RECT 457.380 51.535 457.660 51.815 ;
        RECT 457.380 50.875 457.660 51.155 ;
        RECT 457.380 50.215 457.660 50.495 ;
        RECT 467.665 58.795 467.945 59.075 ;
        RECT 469.085 58.795 469.365 59.075 ;
        RECT 467.665 58.135 467.945 58.415 ;
        RECT 469.085 58.135 469.365 58.415 ;
        RECT 467.665 57.475 467.945 57.755 ;
        RECT 469.085 57.475 469.365 57.755 ;
        RECT 467.665 56.815 467.945 57.095 ;
        RECT 469.085 56.815 469.365 57.095 ;
        RECT 467.665 56.155 467.945 56.435 ;
        RECT 469.085 56.155 469.365 56.435 ;
        RECT 467.665 55.495 467.945 55.775 ;
        RECT 469.085 55.495 469.365 55.775 ;
        RECT 467.665 54.835 467.945 55.115 ;
        RECT 469.085 54.835 469.365 55.115 ;
        RECT 467.665 54.175 467.945 54.455 ;
        RECT 469.085 54.175 469.365 54.455 ;
        RECT 467.665 53.515 467.945 53.795 ;
        RECT 469.085 53.515 469.365 53.795 ;
        RECT 467.665 52.855 467.945 53.135 ;
        RECT 469.085 52.855 469.365 53.135 ;
        RECT 467.665 52.195 467.945 52.475 ;
        RECT 469.085 52.195 469.365 52.475 ;
        RECT 467.665 51.535 467.945 51.815 ;
        RECT 469.085 51.535 469.365 51.815 ;
        RECT 467.665 50.875 467.945 51.155 ;
        RECT 469.085 50.875 469.365 51.155 ;
        RECT 467.665 50.215 467.945 50.495 ;
        RECT 469.085 50.215 469.365 50.495 ;
        RECT 473.570 47.855 473.850 48.135 ;
        RECT 474.230 47.855 474.510 48.135 ;
        RECT 474.890 47.855 475.170 48.135 ;
        RECT 473.570 47.195 473.850 47.475 ;
        RECT 474.230 47.195 474.510 47.475 ;
        RECT 474.890 47.195 475.170 47.475 ;
        RECT 473.570 46.535 473.850 46.815 ;
        RECT 474.230 46.535 474.510 46.815 ;
        RECT 474.890 46.535 475.170 46.815 ;
        RECT 461.875 39.755 462.155 40.035 ;
        RECT 462.535 39.755 462.815 40.035 ;
        RECT 463.195 39.755 463.475 40.035 ;
        RECT 461.875 39.095 462.155 39.375 ;
        RECT 462.535 39.095 462.815 39.375 ;
        RECT 463.195 39.095 463.475 39.375 ;
        RECT 461.875 38.435 462.155 38.715 ;
        RECT 462.535 38.435 462.815 38.715 ;
        RECT 463.195 38.435 463.475 38.715 ;
        RECT 461.875 30.355 462.155 30.635 ;
        RECT 462.535 30.355 462.815 30.635 ;
        RECT 463.195 30.355 463.475 30.635 ;
        RECT 461.875 29.695 462.155 29.975 ;
        RECT 462.535 29.695 462.815 29.975 ;
        RECT 463.195 29.695 463.475 29.975 ;
        RECT 461.875 29.035 462.155 29.315 ;
        RECT 462.535 29.035 462.815 29.315 ;
        RECT 463.195 29.035 463.475 29.315 ;
        RECT 473.570 22.255 473.850 22.535 ;
        RECT 474.230 22.255 474.510 22.535 ;
        RECT 474.890 22.255 475.170 22.535 ;
        RECT 473.570 21.595 473.850 21.875 ;
        RECT 474.230 21.595 474.510 21.875 ;
        RECT 474.890 21.595 475.170 21.875 ;
        RECT 473.570 20.935 473.850 21.215 ;
        RECT 474.230 20.935 474.510 21.215 ;
        RECT 474.890 20.935 475.170 21.215 ;
        RECT 399.440 4.740 399.720 5.020 ;
        RECT 400.100 4.740 400.380 5.020 ;
        RECT 400.760 4.740 401.040 5.020 ;
        RECT 401.680 4.740 401.960 5.020 ;
        RECT 402.340 4.740 402.620 5.020 ;
        RECT 403.000 4.740 403.280 5.020 ;
        RECT 404.040 4.740 404.320 5.020 ;
        RECT 405.040 4.740 405.320 5.020 ;
        RECT 405.700 4.740 405.980 5.020 ;
        RECT 406.360 4.740 406.640 5.020 ;
        RECT 407.280 4.740 407.560 5.020 ;
        RECT 407.940 4.740 408.220 5.020 ;
        RECT 408.600 4.740 408.880 5.020 ;
        RECT 409.520 4.740 409.800 5.020 ;
        RECT 410.180 4.740 410.460 5.020 ;
        RECT 410.840 4.740 411.120 5.020 ;
        RECT 411.760 4.740 412.040 5.020 ;
        RECT 412.420 4.740 412.700 5.020 ;
        RECT 413.080 4.740 413.360 5.020 ;
        RECT 414.000 4.740 414.280 5.020 ;
        RECT 414.660 4.740 414.940 5.020 ;
        RECT 415.320 4.740 415.600 5.020 ;
        RECT 416.240 4.740 416.520 5.020 ;
        RECT 416.900 4.740 417.180 5.020 ;
        RECT 417.560 4.740 417.840 5.020 ;
        RECT 418.480 4.740 418.760 5.020 ;
        RECT 419.140 4.740 419.420 5.020 ;
        RECT 419.800 4.740 420.080 5.020 ;
        RECT 420.720 4.740 421.000 5.020 ;
        RECT 421.380 4.740 421.660 5.020 ;
        RECT 422.040 4.740 422.320 5.020 ;
        RECT 422.960 4.740 423.240 5.020 ;
        RECT 423.620 4.740 423.900 5.020 ;
        RECT 424.280 4.740 424.560 5.020 ;
        RECT 425.320 4.740 425.600 5.020 ;
        RECT 426.320 4.740 426.600 5.020 ;
        RECT 426.980 4.740 427.260 5.020 ;
        RECT 427.640 4.740 427.920 5.020 ;
        RECT 428.560 4.740 428.840 5.020 ;
        RECT 429.220 4.740 429.500 5.020 ;
        RECT 429.880 4.740 430.160 5.020 ;
        RECT 430.800 4.740 431.080 5.020 ;
        RECT 431.460 4.740 431.740 5.020 ;
        RECT 432.120 4.740 432.400 5.020 ;
        RECT 433.040 4.740 433.320 5.020 ;
        RECT 433.700 4.740 433.980 5.020 ;
        RECT 434.360 4.740 434.640 5.020 ;
        RECT 435.280 4.740 435.560 5.020 ;
        RECT 435.940 4.740 436.220 5.020 ;
        RECT 436.600 4.740 436.880 5.020 ;
        RECT 437.620 4.740 437.900 5.020 ;
        RECT 438.280 4.740 438.560 5.020 ;
        RECT 438.940 4.740 439.220 5.020 ;
        RECT 479.375 58.795 479.655 59.075 ;
        RECT 479.375 58.135 479.655 58.415 ;
        RECT 479.375 57.475 479.655 57.755 ;
        RECT 479.375 56.815 479.655 57.095 ;
        RECT 479.375 56.155 479.655 56.435 ;
        RECT 479.375 55.495 479.655 55.775 ;
        RECT 479.375 54.835 479.655 55.115 ;
        RECT 479.375 54.175 479.655 54.455 ;
        RECT 479.375 53.515 479.655 53.795 ;
        RECT 479.375 52.855 479.655 53.135 ;
        RECT 479.375 52.195 479.655 52.475 ;
        RECT 479.375 51.535 479.655 51.815 ;
        RECT 479.375 50.875 479.655 51.155 ;
        RECT 479.375 50.215 479.655 50.495 ;
        RECT 489.660 58.795 489.940 59.075 ;
        RECT 489.660 58.135 489.940 58.415 ;
        RECT 489.660 57.475 489.940 57.755 ;
        RECT 489.660 56.815 489.940 57.095 ;
        RECT 489.660 56.155 489.940 56.435 ;
        RECT 489.660 55.495 489.940 55.775 ;
        RECT 489.660 54.835 489.940 55.115 ;
        RECT 489.660 54.175 489.940 54.455 ;
        RECT 489.660 53.515 489.940 53.795 ;
        RECT 489.660 52.855 489.940 53.135 ;
        RECT 489.660 52.195 489.940 52.475 ;
        RECT 489.660 51.535 489.940 51.815 ;
        RECT 489.660 50.875 489.940 51.155 ;
        RECT 489.660 50.215 489.940 50.495 ;
        RECT 483.870 45.155 484.150 45.435 ;
        RECT 484.530 45.155 484.810 45.435 ;
        RECT 485.190 45.155 485.470 45.435 ;
        RECT 483.870 44.495 484.150 44.775 ;
        RECT 484.530 44.495 484.810 44.775 ;
        RECT 485.190 44.495 485.470 44.775 ;
        RECT 483.870 43.835 484.150 44.115 ;
        RECT 484.530 43.835 484.810 44.115 ;
        RECT 485.190 43.835 485.470 44.115 ;
        RECT 494.145 42.455 494.425 42.735 ;
        RECT 494.805 42.455 495.085 42.735 ;
        RECT 495.465 42.455 495.745 42.735 ;
        RECT 494.145 41.795 494.425 42.075 ;
        RECT 494.805 41.795 495.085 42.075 ;
        RECT 495.465 41.795 495.745 42.075 ;
        RECT 494.145 41.135 494.425 41.415 ;
        RECT 494.805 41.135 495.085 41.415 ;
        RECT 495.465 41.135 495.745 41.415 ;
        RECT 494.145 27.655 494.425 27.935 ;
        RECT 494.805 27.655 495.085 27.935 ;
        RECT 495.465 27.655 495.745 27.935 ;
        RECT 494.145 26.995 494.425 27.275 ;
        RECT 494.805 26.995 495.085 27.275 ;
        RECT 495.465 26.995 495.745 27.275 ;
        RECT 494.145 26.335 494.425 26.615 ;
        RECT 494.805 26.335 495.085 26.615 ;
        RECT 495.465 26.335 495.745 26.615 ;
        RECT 483.870 24.955 484.150 25.235 ;
        RECT 484.530 24.955 484.810 25.235 ;
        RECT 485.190 24.955 485.470 25.235 ;
        RECT 483.870 24.295 484.150 24.575 ;
        RECT 484.530 24.295 484.810 24.575 ;
        RECT 485.190 24.295 485.470 24.575 ;
        RECT 483.870 23.635 484.150 23.915 ;
        RECT 484.530 23.635 484.810 23.915 ;
        RECT 485.190 23.635 485.470 23.915 ;
        RECT 499.950 58.795 500.230 59.075 ;
        RECT 499.950 58.135 500.230 58.415 ;
        RECT 499.950 57.475 500.230 57.755 ;
        RECT 499.950 56.815 500.230 57.095 ;
        RECT 499.950 56.155 500.230 56.435 ;
        RECT 499.950 55.495 500.230 55.775 ;
        RECT 499.950 54.835 500.230 55.115 ;
        RECT 499.950 54.175 500.230 54.455 ;
        RECT 499.950 53.515 500.230 53.795 ;
        RECT 499.950 52.855 500.230 53.135 ;
        RECT 499.950 52.195 500.230 52.475 ;
        RECT 499.950 51.535 500.230 51.815 ;
        RECT 499.950 50.875 500.230 51.155 ;
        RECT 499.950 50.215 500.230 50.495 ;
        RECT 510.235 58.795 510.515 59.075 ;
        RECT 511.655 58.795 511.935 59.075 ;
        RECT 510.235 58.135 510.515 58.415 ;
        RECT 511.655 58.135 511.935 58.415 ;
        RECT 510.235 57.475 510.515 57.755 ;
        RECT 511.655 57.475 511.935 57.755 ;
        RECT 510.235 56.815 510.515 57.095 ;
        RECT 511.655 56.815 511.935 57.095 ;
        RECT 510.235 56.155 510.515 56.435 ;
        RECT 511.655 56.155 511.935 56.435 ;
        RECT 510.235 55.495 510.515 55.775 ;
        RECT 511.655 55.495 511.935 55.775 ;
        RECT 510.235 54.835 510.515 55.115 ;
        RECT 511.655 54.835 511.935 55.115 ;
        RECT 510.235 54.175 510.515 54.455 ;
        RECT 511.655 54.175 511.935 54.455 ;
        RECT 510.235 53.515 510.515 53.795 ;
        RECT 511.655 53.515 511.935 53.795 ;
        RECT 510.235 52.855 510.515 53.135 ;
        RECT 511.655 52.855 511.935 53.135 ;
        RECT 510.235 52.195 510.515 52.475 ;
        RECT 511.655 52.195 511.935 52.475 ;
        RECT 510.235 51.535 510.515 51.815 ;
        RECT 511.655 51.535 511.935 51.815 ;
        RECT 510.235 50.875 510.515 51.155 ;
        RECT 511.655 50.875 511.935 51.155 ;
        RECT 510.235 50.215 510.515 50.495 ;
        RECT 511.655 50.215 511.935 50.495 ;
        RECT 516.140 47.855 516.420 48.135 ;
        RECT 516.800 47.855 517.080 48.135 ;
        RECT 517.460 47.855 517.740 48.135 ;
        RECT 516.140 47.195 516.420 47.475 ;
        RECT 516.800 47.195 517.080 47.475 ;
        RECT 517.460 47.195 517.740 47.475 ;
        RECT 516.140 46.535 516.420 46.815 ;
        RECT 516.800 46.535 517.080 46.815 ;
        RECT 517.460 46.535 517.740 46.815 ;
        RECT 504.445 39.755 504.725 40.035 ;
        RECT 505.105 39.755 505.385 40.035 ;
        RECT 505.765 39.755 506.045 40.035 ;
        RECT 504.445 39.095 504.725 39.375 ;
        RECT 505.105 39.095 505.385 39.375 ;
        RECT 505.765 39.095 506.045 39.375 ;
        RECT 504.445 38.435 504.725 38.715 ;
        RECT 505.105 38.435 505.385 38.715 ;
        RECT 505.765 38.435 506.045 38.715 ;
        RECT 504.445 30.355 504.725 30.635 ;
        RECT 505.105 30.355 505.385 30.635 ;
        RECT 505.765 30.355 506.045 30.635 ;
        RECT 504.445 29.695 504.725 29.975 ;
        RECT 505.105 29.695 505.385 29.975 ;
        RECT 505.765 29.695 506.045 29.975 ;
        RECT 504.445 29.035 504.725 29.315 ;
        RECT 505.105 29.035 505.385 29.315 ;
        RECT 505.765 29.035 506.045 29.315 ;
        RECT 516.140 22.255 516.420 22.535 ;
        RECT 516.800 22.255 517.080 22.535 ;
        RECT 517.460 22.255 517.740 22.535 ;
        RECT 516.140 21.595 516.420 21.875 ;
        RECT 516.800 21.595 517.080 21.875 ;
        RECT 517.460 21.595 517.740 21.875 ;
        RECT 516.140 20.935 516.420 21.215 ;
        RECT 516.800 20.935 517.080 21.215 ;
        RECT 517.460 20.935 517.740 21.215 ;
        RECT 440.880 4.740 441.160 5.020 ;
        RECT 441.540 4.740 441.820 5.020 ;
        RECT 442.200 4.740 442.480 5.020 ;
        RECT 443.120 4.740 443.400 5.020 ;
        RECT 443.780 4.740 444.060 5.020 ;
        RECT 444.440 4.740 444.720 5.020 ;
        RECT 445.480 4.740 445.760 5.020 ;
        RECT 446.480 4.740 446.760 5.020 ;
        RECT 447.140 4.740 447.420 5.020 ;
        RECT 447.800 4.740 448.080 5.020 ;
        RECT 448.720 4.740 449.000 5.020 ;
        RECT 449.380 4.740 449.660 5.020 ;
        RECT 450.040 4.740 450.320 5.020 ;
        RECT 450.960 4.740 451.240 5.020 ;
        RECT 451.620 4.740 451.900 5.020 ;
        RECT 452.280 4.740 452.560 5.020 ;
        RECT 453.200 4.740 453.480 5.020 ;
        RECT 453.860 4.740 454.140 5.020 ;
        RECT 454.520 4.740 454.800 5.020 ;
        RECT 455.440 4.740 455.720 5.020 ;
        RECT 456.100 4.740 456.380 5.020 ;
        RECT 456.760 4.740 457.040 5.020 ;
        RECT 457.680 4.740 457.960 5.020 ;
        RECT 458.340 4.740 458.620 5.020 ;
        RECT 459.000 4.740 459.280 5.020 ;
        RECT 459.920 4.740 460.200 5.020 ;
        RECT 460.580 4.740 460.860 5.020 ;
        RECT 461.240 4.740 461.520 5.020 ;
        RECT 462.160 4.740 462.440 5.020 ;
        RECT 462.820 4.740 463.100 5.020 ;
        RECT 463.480 4.740 463.760 5.020 ;
        RECT 464.400 4.740 464.680 5.020 ;
        RECT 465.060 4.740 465.340 5.020 ;
        RECT 465.720 4.740 466.000 5.020 ;
        RECT 466.760 4.740 467.040 5.020 ;
        RECT 467.760 4.740 468.040 5.020 ;
        RECT 468.420 4.740 468.700 5.020 ;
        RECT 469.080 4.740 469.360 5.020 ;
        RECT 470.000 4.740 470.280 5.020 ;
        RECT 470.660 4.740 470.940 5.020 ;
        RECT 471.320 4.740 471.600 5.020 ;
        RECT 472.240 4.740 472.520 5.020 ;
        RECT 472.900 4.740 473.180 5.020 ;
        RECT 473.560 4.740 473.840 5.020 ;
        RECT 474.480 4.740 474.760 5.020 ;
        RECT 475.140 4.740 475.420 5.020 ;
        RECT 475.800 4.740 476.080 5.020 ;
        RECT 476.720 4.740 477.000 5.020 ;
        RECT 477.380 4.740 477.660 5.020 ;
        RECT 478.040 4.740 478.320 5.020 ;
        RECT 478.960 4.740 479.240 5.020 ;
        RECT 479.620 4.740 479.900 5.020 ;
        RECT 480.280 4.740 480.560 5.020 ;
        RECT 481.300 4.740 481.580 5.020 ;
        RECT 481.960 4.740 482.240 5.020 ;
        RECT 482.620 4.740 482.900 5.020 ;
        RECT 521.945 58.795 522.225 59.075 ;
        RECT 521.945 58.135 522.225 58.415 ;
        RECT 521.945 57.475 522.225 57.755 ;
        RECT 521.945 56.815 522.225 57.095 ;
        RECT 521.945 56.155 522.225 56.435 ;
        RECT 521.945 55.495 522.225 55.775 ;
        RECT 521.945 54.835 522.225 55.115 ;
        RECT 521.945 54.175 522.225 54.455 ;
        RECT 521.945 53.515 522.225 53.795 ;
        RECT 521.945 52.855 522.225 53.135 ;
        RECT 521.945 52.195 522.225 52.475 ;
        RECT 521.945 51.535 522.225 51.815 ;
        RECT 521.945 50.875 522.225 51.155 ;
        RECT 521.945 50.215 522.225 50.495 ;
        RECT 532.230 58.795 532.510 59.075 ;
        RECT 532.230 58.135 532.510 58.415 ;
        RECT 532.230 57.475 532.510 57.755 ;
        RECT 532.230 56.815 532.510 57.095 ;
        RECT 532.230 56.155 532.510 56.435 ;
        RECT 532.230 55.495 532.510 55.775 ;
        RECT 532.230 54.835 532.510 55.115 ;
        RECT 532.230 54.175 532.510 54.455 ;
        RECT 532.230 53.515 532.510 53.795 ;
        RECT 532.230 52.855 532.510 53.135 ;
        RECT 532.230 52.195 532.510 52.475 ;
        RECT 532.230 51.535 532.510 51.815 ;
        RECT 532.230 50.875 532.510 51.155 ;
        RECT 532.230 50.215 532.510 50.495 ;
        RECT 526.440 45.155 526.720 45.435 ;
        RECT 527.100 45.155 527.380 45.435 ;
        RECT 527.760 45.155 528.040 45.435 ;
        RECT 526.440 44.495 526.720 44.775 ;
        RECT 527.100 44.495 527.380 44.775 ;
        RECT 527.760 44.495 528.040 44.775 ;
        RECT 526.440 43.835 526.720 44.115 ;
        RECT 527.100 43.835 527.380 44.115 ;
        RECT 527.760 43.835 528.040 44.115 ;
        RECT 536.715 42.455 536.995 42.735 ;
        RECT 537.375 42.455 537.655 42.735 ;
        RECT 538.035 42.455 538.315 42.735 ;
        RECT 536.715 41.795 536.995 42.075 ;
        RECT 537.375 41.795 537.655 42.075 ;
        RECT 538.035 41.795 538.315 42.075 ;
        RECT 536.715 41.135 536.995 41.415 ;
        RECT 537.375 41.135 537.655 41.415 ;
        RECT 538.035 41.135 538.315 41.415 ;
        RECT 536.715 27.655 536.995 27.935 ;
        RECT 537.375 27.655 537.655 27.935 ;
        RECT 538.035 27.655 538.315 27.935 ;
        RECT 536.715 26.995 536.995 27.275 ;
        RECT 537.375 26.995 537.655 27.275 ;
        RECT 538.035 26.995 538.315 27.275 ;
        RECT 536.715 26.335 536.995 26.615 ;
        RECT 537.375 26.335 537.655 26.615 ;
        RECT 538.035 26.335 538.315 26.615 ;
        RECT 526.440 24.955 526.720 25.235 ;
        RECT 527.100 24.955 527.380 25.235 ;
        RECT 527.760 24.955 528.040 25.235 ;
        RECT 526.440 24.295 526.720 24.575 ;
        RECT 527.100 24.295 527.380 24.575 ;
        RECT 527.760 24.295 528.040 24.575 ;
        RECT 526.440 23.635 526.720 23.915 ;
        RECT 527.100 23.635 527.380 23.915 ;
        RECT 527.760 23.635 528.040 23.915 ;
        RECT 542.520 58.795 542.800 59.075 ;
        RECT 542.520 58.135 542.800 58.415 ;
        RECT 542.520 57.475 542.800 57.755 ;
        RECT 542.520 56.815 542.800 57.095 ;
        RECT 542.520 56.155 542.800 56.435 ;
        RECT 542.520 55.495 542.800 55.775 ;
        RECT 542.520 54.835 542.800 55.115 ;
        RECT 542.520 54.175 542.800 54.455 ;
        RECT 542.520 53.515 542.800 53.795 ;
        RECT 542.520 52.855 542.800 53.135 ;
        RECT 542.520 52.195 542.800 52.475 ;
        RECT 542.520 51.535 542.800 51.815 ;
        RECT 542.520 50.875 542.800 51.155 ;
        RECT 542.520 50.215 542.800 50.495 ;
        RECT 552.805 58.795 553.085 59.075 ;
        RECT 554.225 58.795 554.505 59.075 ;
        RECT 552.805 58.135 553.085 58.415 ;
        RECT 554.225 58.135 554.505 58.415 ;
        RECT 552.805 57.475 553.085 57.755 ;
        RECT 554.225 57.475 554.505 57.755 ;
        RECT 552.805 56.815 553.085 57.095 ;
        RECT 554.225 56.815 554.505 57.095 ;
        RECT 552.805 56.155 553.085 56.435 ;
        RECT 554.225 56.155 554.505 56.435 ;
        RECT 552.805 55.495 553.085 55.775 ;
        RECT 554.225 55.495 554.505 55.775 ;
        RECT 552.805 54.835 553.085 55.115 ;
        RECT 554.225 54.835 554.505 55.115 ;
        RECT 552.805 54.175 553.085 54.455 ;
        RECT 554.225 54.175 554.505 54.455 ;
        RECT 552.805 53.515 553.085 53.795 ;
        RECT 554.225 53.515 554.505 53.795 ;
        RECT 552.805 52.855 553.085 53.135 ;
        RECT 554.225 52.855 554.505 53.135 ;
        RECT 552.805 52.195 553.085 52.475 ;
        RECT 554.225 52.195 554.505 52.475 ;
        RECT 552.805 51.535 553.085 51.815 ;
        RECT 554.225 51.535 554.505 51.815 ;
        RECT 552.805 50.875 553.085 51.155 ;
        RECT 554.225 50.875 554.505 51.155 ;
        RECT 552.805 50.215 553.085 50.495 ;
        RECT 554.225 50.215 554.505 50.495 ;
        RECT 558.710 47.855 558.990 48.135 ;
        RECT 559.370 47.855 559.650 48.135 ;
        RECT 560.030 47.855 560.310 48.135 ;
        RECT 558.710 47.195 558.990 47.475 ;
        RECT 559.370 47.195 559.650 47.475 ;
        RECT 560.030 47.195 560.310 47.475 ;
        RECT 558.710 46.535 558.990 46.815 ;
        RECT 559.370 46.535 559.650 46.815 ;
        RECT 560.030 46.535 560.310 46.815 ;
        RECT 547.015 39.755 547.295 40.035 ;
        RECT 547.675 39.755 547.955 40.035 ;
        RECT 548.335 39.755 548.615 40.035 ;
        RECT 547.015 39.095 547.295 39.375 ;
        RECT 547.675 39.095 547.955 39.375 ;
        RECT 548.335 39.095 548.615 39.375 ;
        RECT 547.015 38.435 547.295 38.715 ;
        RECT 547.675 38.435 547.955 38.715 ;
        RECT 548.335 38.435 548.615 38.715 ;
        RECT 547.015 30.355 547.295 30.635 ;
        RECT 547.675 30.355 547.955 30.635 ;
        RECT 548.335 30.355 548.615 30.635 ;
        RECT 547.015 29.695 547.295 29.975 ;
        RECT 547.675 29.695 547.955 29.975 ;
        RECT 548.335 29.695 548.615 29.975 ;
        RECT 547.015 29.035 547.295 29.315 ;
        RECT 547.675 29.035 547.955 29.315 ;
        RECT 548.335 29.035 548.615 29.315 ;
        RECT 558.710 22.255 558.990 22.535 ;
        RECT 559.370 22.255 559.650 22.535 ;
        RECT 560.030 22.255 560.310 22.535 ;
        RECT 558.710 21.595 558.990 21.875 ;
        RECT 559.370 21.595 559.650 21.875 ;
        RECT 560.030 21.595 560.310 21.875 ;
        RECT 558.710 20.935 558.990 21.215 ;
        RECT 559.370 20.935 559.650 21.215 ;
        RECT 560.030 20.935 560.310 21.215 ;
        RECT 484.560 4.740 484.840 5.020 ;
        RECT 485.220 4.740 485.500 5.020 ;
        RECT 485.880 4.740 486.160 5.020 ;
        RECT 486.920 4.740 487.200 5.020 ;
        RECT 487.920 4.740 488.200 5.020 ;
        RECT 488.580 4.740 488.860 5.020 ;
        RECT 489.240 4.740 489.520 5.020 ;
        RECT 490.160 4.740 490.440 5.020 ;
        RECT 490.820 4.740 491.100 5.020 ;
        RECT 491.480 4.740 491.760 5.020 ;
        RECT 492.400 4.740 492.680 5.020 ;
        RECT 493.060 4.740 493.340 5.020 ;
        RECT 493.720 4.740 494.000 5.020 ;
        RECT 494.640 4.740 494.920 5.020 ;
        RECT 495.300 4.740 495.580 5.020 ;
        RECT 495.960 4.740 496.240 5.020 ;
        RECT 496.880 4.740 497.160 5.020 ;
        RECT 497.540 4.740 497.820 5.020 ;
        RECT 498.200 4.740 498.480 5.020 ;
        RECT 499.120 4.740 499.400 5.020 ;
        RECT 499.780 4.740 500.060 5.020 ;
        RECT 500.440 4.740 500.720 5.020 ;
        RECT 501.360 4.740 501.640 5.020 ;
        RECT 502.020 4.740 502.300 5.020 ;
        RECT 502.680 4.740 502.960 5.020 ;
        RECT 503.600 4.740 503.880 5.020 ;
        RECT 504.260 4.740 504.540 5.020 ;
        RECT 504.920 4.740 505.200 5.020 ;
        RECT 505.840 4.740 506.120 5.020 ;
        RECT 506.500 4.740 506.780 5.020 ;
        RECT 507.160 4.740 507.440 5.020 ;
        RECT 508.200 4.740 508.480 5.020 ;
        RECT 509.200 4.740 509.480 5.020 ;
        RECT 509.860 4.740 510.140 5.020 ;
        RECT 510.520 4.740 510.800 5.020 ;
        RECT 511.440 4.740 511.720 5.020 ;
        RECT 512.100 4.740 512.380 5.020 ;
        RECT 512.760 4.740 513.040 5.020 ;
        RECT 513.680 4.740 513.960 5.020 ;
        RECT 514.340 4.740 514.620 5.020 ;
        RECT 515.000 4.740 515.280 5.020 ;
        RECT 515.920 4.740 516.200 5.020 ;
        RECT 516.580 4.740 516.860 5.020 ;
        RECT 517.240 4.740 517.520 5.020 ;
        RECT 518.160 4.740 518.440 5.020 ;
        RECT 518.820 4.740 519.100 5.020 ;
        RECT 519.480 4.740 519.760 5.020 ;
        RECT 520.400 4.740 520.680 5.020 ;
        RECT 521.060 4.740 521.340 5.020 ;
        RECT 521.720 4.740 522.000 5.020 ;
        RECT 522.740 4.740 523.020 5.020 ;
        RECT 523.400 4.740 523.680 5.020 ;
        RECT 524.060 4.740 524.340 5.020 ;
        RECT 564.515 58.795 564.795 59.075 ;
        RECT 564.515 58.135 564.795 58.415 ;
        RECT 564.515 57.475 564.795 57.755 ;
        RECT 564.515 56.815 564.795 57.095 ;
        RECT 564.515 56.155 564.795 56.435 ;
        RECT 564.515 55.495 564.795 55.775 ;
        RECT 564.515 54.835 564.795 55.115 ;
        RECT 564.515 54.175 564.795 54.455 ;
        RECT 564.515 53.515 564.795 53.795 ;
        RECT 564.515 52.855 564.795 53.135 ;
        RECT 564.515 52.195 564.795 52.475 ;
        RECT 564.515 51.535 564.795 51.815 ;
        RECT 564.515 50.875 564.795 51.155 ;
        RECT 564.515 50.215 564.795 50.495 ;
        RECT 574.800 58.795 575.080 59.075 ;
        RECT 574.800 58.135 575.080 58.415 ;
        RECT 574.800 57.475 575.080 57.755 ;
        RECT 574.800 56.815 575.080 57.095 ;
        RECT 574.800 56.155 575.080 56.435 ;
        RECT 574.800 55.495 575.080 55.775 ;
        RECT 574.800 54.835 575.080 55.115 ;
        RECT 574.800 54.175 575.080 54.455 ;
        RECT 574.800 53.515 575.080 53.795 ;
        RECT 574.800 52.855 575.080 53.135 ;
        RECT 574.800 52.195 575.080 52.475 ;
        RECT 574.800 51.535 575.080 51.815 ;
        RECT 574.800 50.875 575.080 51.155 ;
        RECT 574.800 50.215 575.080 50.495 ;
        RECT 569.010 45.155 569.290 45.435 ;
        RECT 569.670 45.155 569.950 45.435 ;
        RECT 570.330 45.155 570.610 45.435 ;
        RECT 569.010 44.495 569.290 44.775 ;
        RECT 569.670 44.495 569.950 44.775 ;
        RECT 570.330 44.495 570.610 44.775 ;
        RECT 569.010 43.835 569.290 44.115 ;
        RECT 569.670 43.835 569.950 44.115 ;
        RECT 570.330 43.835 570.610 44.115 ;
        RECT 579.285 42.455 579.565 42.735 ;
        RECT 579.945 42.455 580.225 42.735 ;
        RECT 580.605 42.455 580.885 42.735 ;
        RECT 579.285 41.795 579.565 42.075 ;
        RECT 579.945 41.795 580.225 42.075 ;
        RECT 580.605 41.795 580.885 42.075 ;
        RECT 579.285 41.135 579.565 41.415 ;
        RECT 579.945 41.135 580.225 41.415 ;
        RECT 580.605 41.135 580.885 41.415 ;
        RECT 579.285 27.655 579.565 27.935 ;
        RECT 579.945 27.655 580.225 27.935 ;
        RECT 580.605 27.655 580.885 27.935 ;
        RECT 579.285 26.995 579.565 27.275 ;
        RECT 579.945 26.995 580.225 27.275 ;
        RECT 580.605 26.995 580.885 27.275 ;
        RECT 579.285 26.335 579.565 26.615 ;
        RECT 579.945 26.335 580.225 26.615 ;
        RECT 580.605 26.335 580.885 26.615 ;
        RECT 569.010 24.955 569.290 25.235 ;
        RECT 569.670 24.955 569.950 25.235 ;
        RECT 570.330 24.955 570.610 25.235 ;
        RECT 569.010 24.295 569.290 24.575 ;
        RECT 569.670 24.295 569.950 24.575 ;
        RECT 570.330 24.295 570.610 24.575 ;
        RECT 569.010 23.635 569.290 23.915 ;
        RECT 569.670 23.635 569.950 23.915 ;
        RECT 570.330 23.635 570.610 23.915 ;
        RECT 585.090 58.795 585.370 59.075 ;
        RECT 585.090 58.135 585.370 58.415 ;
        RECT 585.090 57.475 585.370 57.755 ;
        RECT 585.090 56.815 585.370 57.095 ;
        RECT 585.090 56.155 585.370 56.435 ;
        RECT 585.090 55.495 585.370 55.775 ;
        RECT 585.090 54.835 585.370 55.115 ;
        RECT 585.090 54.175 585.370 54.455 ;
        RECT 585.090 53.515 585.370 53.795 ;
        RECT 585.090 52.855 585.370 53.135 ;
        RECT 585.090 52.195 585.370 52.475 ;
        RECT 585.090 51.535 585.370 51.815 ;
        RECT 585.090 50.875 585.370 51.155 ;
        RECT 585.090 50.215 585.370 50.495 ;
        RECT 595.375 58.795 595.655 59.075 ;
        RECT 596.795 58.795 597.075 59.075 ;
        RECT 595.375 58.135 595.655 58.415 ;
        RECT 596.795 58.135 597.075 58.415 ;
        RECT 595.375 57.475 595.655 57.755 ;
        RECT 596.795 57.475 597.075 57.755 ;
        RECT 595.375 56.815 595.655 57.095 ;
        RECT 596.795 56.815 597.075 57.095 ;
        RECT 595.375 56.155 595.655 56.435 ;
        RECT 596.795 56.155 597.075 56.435 ;
        RECT 595.375 55.495 595.655 55.775 ;
        RECT 596.795 55.495 597.075 55.775 ;
        RECT 595.375 54.835 595.655 55.115 ;
        RECT 596.795 54.835 597.075 55.115 ;
        RECT 595.375 54.175 595.655 54.455 ;
        RECT 596.795 54.175 597.075 54.455 ;
        RECT 595.375 53.515 595.655 53.795 ;
        RECT 596.795 53.515 597.075 53.795 ;
        RECT 595.375 52.855 595.655 53.135 ;
        RECT 596.795 52.855 597.075 53.135 ;
        RECT 595.375 52.195 595.655 52.475 ;
        RECT 596.795 52.195 597.075 52.475 ;
        RECT 595.375 51.535 595.655 51.815 ;
        RECT 596.795 51.535 597.075 51.815 ;
        RECT 595.375 50.875 595.655 51.155 ;
        RECT 596.795 50.875 597.075 51.155 ;
        RECT 595.375 50.215 595.655 50.495 ;
        RECT 596.795 50.215 597.075 50.495 ;
        RECT 601.280 47.855 601.560 48.135 ;
        RECT 601.940 47.855 602.220 48.135 ;
        RECT 602.600 47.855 602.880 48.135 ;
        RECT 601.280 47.195 601.560 47.475 ;
        RECT 601.940 47.195 602.220 47.475 ;
        RECT 602.600 47.195 602.880 47.475 ;
        RECT 601.280 46.535 601.560 46.815 ;
        RECT 601.940 46.535 602.220 46.815 ;
        RECT 602.600 46.535 602.880 46.815 ;
        RECT 589.585 39.755 589.865 40.035 ;
        RECT 590.245 39.755 590.525 40.035 ;
        RECT 590.905 39.755 591.185 40.035 ;
        RECT 589.585 39.095 589.865 39.375 ;
        RECT 590.245 39.095 590.525 39.375 ;
        RECT 590.905 39.095 591.185 39.375 ;
        RECT 589.585 38.435 589.865 38.715 ;
        RECT 590.245 38.435 590.525 38.715 ;
        RECT 590.905 38.435 591.185 38.715 ;
        RECT 589.585 30.355 589.865 30.635 ;
        RECT 590.245 30.355 590.525 30.635 ;
        RECT 590.905 30.355 591.185 30.635 ;
        RECT 589.585 29.695 589.865 29.975 ;
        RECT 590.245 29.695 590.525 29.975 ;
        RECT 590.905 29.695 591.185 29.975 ;
        RECT 589.585 29.035 589.865 29.315 ;
        RECT 590.245 29.035 590.525 29.315 ;
        RECT 590.905 29.035 591.185 29.315 ;
        RECT 601.280 22.255 601.560 22.535 ;
        RECT 601.940 22.255 602.220 22.535 ;
        RECT 602.600 22.255 602.880 22.535 ;
        RECT 601.280 21.595 601.560 21.875 ;
        RECT 601.940 21.595 602.220 21.875 ;
        RECT 602.600 21.595 602.880 21.875 ;
        RECT 601.280 20.935 601.560 21.215 ;
        RECT 601.940 20.935 602.220 21.215 ;
        RECT 602.600 20.935 602.880 21.215 ;
        RECT 526.000 4.740 526.280 5.020 ;
        RECT 526.660 4.740 526.940 5.020 ;
        RECT 527.320 4.740 527.600 5.020 ;
        RECT 528.360 4.740 528.640 5.020 ;
        RECT 529.360 4.740 529.640 5.020 ;
        RECT 530.020 4.740 530.300 5.020 ;
        RECT 530.680 4.740 530.960 5.020 ;
        RECT 531.600 4.740 531.880 5.020 ;
        RECT 532.260 4.740 532.540 5.020 ;
        RECT 532.920 4.740 533.200 5.020 ;
        RECT 533.840 4.740 534.120 5.020 ;
        RECT 534.500 4.740 534.780 5.020 ;
        RECT 535.160 4.740 535.440 5.020 ;
        RECT 536.080 4.740 536.360 5.020 ;
        RECT 536.740 4.740 537.020 5.020 ;
        RECT 537.400 4.740 537.680 5.020 ;
        RECT 538.320 4.740 538.600 5.020 ;
        RECT 538.980 4.740 539.260 5.020 ;
        RECT 539.640 4.740 539.920 5.020 ;
        RECT 540.560 4.740 540.840 5.020 ;
        RECT 541.220 4.740 541.500 5.020 ;
        RECT 541.880 4.740 542.160 5.020 ;
        RECT 542.800 4.740 543.080 5.020 ;
        RECT 543.460 4.740 543.740 5.020 ;
        RECT 544.120 4.740 544.400 5.020 ;
        RECT 545.040 4.740 545.320 5.020 ;
        RECT 545.700 4.740 545.980 5.020 ;
        RECT 546.360 4.740 546.640 5.020 ;
        RECT 547.280 4.740 547.560 5.020 ;
        RECT 547.940 4.740 548.220 5.020 ;
        RECT 548.600 4.740 548.880 5.020 ;
        RECT 549.640 4.740 549.920 5.020 ;
        RECT 550.640 4.740 550.920 5.020 ;
        RECT 551.300 4.740 551.580 5.020 ;
        RECT 551.960 4.740 552.240 5.020 ;
        RECT 552.880 4.740 553.160 5.020 ;
        RECT 553.540 4.740 553.820 5.020 ;
        RECT 554.200 4.740 554.480 5.020 ;
        RECT 555.120 4.740 555.400 5.020 ;
        RECT 555.780 4.740 556.060 5.020 ;
        RECT 556.440 4.740 556.720 5.020 ;
        RECT 557.360 4.740 557.640 5.020 ;
        RECT 558.020 4.740 558.300 5.020 ;
        RECT 558.680 4.740 558.960 5.020 ;
        RECT 559.600 4.740 559.880 5.020 ;
        RECT 560.260 4.740 560.540 5.020 ;
        RECT 560.920 4.740 561.200 5.020 ;
        RECT 561.840 4.740 562.120 5.020 ;
        RECT 562.500 4.740 562.780 5.020 ;
        RECT 563.160 4.740 563.440 5.020 ;
        RECT 564.080 4.740 564.360 5.020 ;
        RECT 564.740 4.740 565.020 5.020 ;
        RECT 565.400 4.740 565.680 5.020 ;
        RECT 566.420 4.740 566.700 5.020 ;
        RECT 567.080 4.740 567.360 5.020 ;
        RECT 567.740 4.740 568.020 5.020 ;
        RECT 607.085 58.795 607.365 59.075 ;
        RECT 607.085 58.135 607.365 58.415 ;
        RECT 607.085 57.475 607.365 57.755 ;
        RECT 607.085 56.815 607.365 57.095 ;
        RECT 607.085 56.155 607.365 56.435 ;
        RECT 607.085 55.495 607.365 55.775 ;
        RECT 607.085 54.835 607.365 55.115 ;
        RECT 607.085 54.175 607.365 54.455 ;
        RECT 607.085 53.515 607.365 53.795 ;
        RECT 607.085 52.855 607.365 53.135 ;
        RECT 607.085 52.195 607.365 52.475 ;
        RECT 607.085 51.535 607.365 51.815 ;
        RECT 607.085 50.875 607.365 51.155 ;
        RECT 607.085 50.215 607.365 50.495 ;
        RECT 617.370 58.795 617.650 59.075 ;
        RECT 617.370 58.135 617.650 58.415 ;
        RECT 617.370 57.475 617.650 57.755 ;
        RECT 617.370 56.815 617.650 57.095 ;
        RECT 617.370 56.155 617.650 56.435 ;
        RECT 617.370 55.495 617.650 55.775 ;
        RECT 617.370 54.835 617.650 55.115 ;
        RECT 617.370 54.175 617.650 54.455 ;
        RECT 617.370 53.515 617.650 53.795 ;
        RECT 617.370 52.855 617.650 53.135 ;
        RECT 617.370 52.195 617.650 52.475 ;
        RECT 617.370 51.535 617.650 51.815 ;
        RECT 617.370 50.875 617.650 51.155 ;
        RECT 617.370 50.215 617.650 50.495 ;
        RECT 611.580 45.155 611.860 45.435 ;
        RECT 612.240 45.155 612.520 45.435 ;
        RECT 612.900 45.155 613.180 45.435 ;
        RECT 611.580 44.495 611.860 44.775 ;
        RECT 612.240 44.495 612.520 44.775 ;
        RECT 612.900 44.495 613.180 44.775 ;
        RECT 611.580 43.835 611.860 44.115 ;
        RECT 612.240 43.835 612.520 44.115 ;
        RECT 612.900 43.835 613.180 44.115 ;
        RECT 621.855 42.455 622.135 42.735 ;
        RECT 622.515 42.455 622.795 42.735 ;
        RECT 623.175 42.455 623.455 42.735 ;
        RECT 621.855 41.795 622.135 42.075 ;
        RECT 622.515 41.795 622.795 42.075 ;
        RECT 623.175 41.795 623.455 42.075 ;
        RECT 621.855 41.135 622.135 41.415 ;
        RECT 622.515 41.135 622.795 41.415 ;
        RECT 623.175 41.135 623.455 41.415 ;
        RECT 621.855 27.655 622.135 27.935 ;
        RECT 622.515 27.655 622.795 27.935 ;
        RECT 623.175 27.655 623.455 27.935 ;
        RECT 621.855 26.995 622.135 27.275 ;
        RECT 622.515 26.995 622.795 27.275 ;
        RECT 623.175 26.995 623.455 27.275 ;
        RECT 621.855 26.335 622.135 26.615 ;
        RECT 622.515 26.335 622.795 26.615 ;
        RECT 623.175 26.335 623.455 26.615 ;
        RECT 611.580 24.955 611.860 25.235 ;
        RECT 612.240 24.955 612.520 25.235 ;
        RECT 612.900 24.955 613.180 25.235 ;
        RECT 611.580 24.295 611.860 24.575 ;
        RECT 612.240 24.295 612.520 24.575 ;
        RECT 612.900 24.295 613.180 24.575 ;
        RECT 611.580 23.635 611.860 23.915 ;
        RECT 612.240 23.635 612.520 23.915 ;
        RECT 612.900 23.635 613.180 23.915 ;
        RECT 627.660 58.795 627.940 59.075 ;
        RECT 627.660 58.135 627.940 58.415 ;
        RECT 627.660 57.475 627.940 57.755 ;
        RECT 627.660 56.815 627.940 57.095 ;
        RECT 627.660 56.155 627.940 56.435 ;
        RECT 627.660 55.495 627.940 55.775 ;
        RECT 627.660 54.835 627.940 55.115 ;
        RECT 627.660 54.175 627.940 54.455 ;
        RECT 627.660 53.515 627.940 53.795 ;
        RECT 627.660 52.855 627.940 53.135 ;
        RECT 627.660 52.195 627.940 52.475 ;
        RECT 627.660 51.535 627.940 51.815 ;
        RECT 627.660 50.875 627.940 51.155 ;
        RECT 627.660 50.215 627.940 50.495 ;
        RECT 637.945 58.795 638.225 59.075 ;
        RECT 639.365 58.795 639.645 59.075 ;
        RECT 637.945 58.135 638.225 58.415 ;
        RECT 639.365 58.135 639.645 58.415 ;
        RECT 637.945 57.475 638.225 57.755 ;
        RECT 639.365 57.475 639.645 57.755 ;
        RECT 637.945 56.815 638.225 57.095 ;
        RECT 639.365 56.815 639.645 57.095 ;
        RECT 637.945 56.155 638.225 56.435 ;
        RECT 639.365 56.155 639.645 56.435 ;
        RECT 637.945 55.495 638.225 55.775 ;
        RECT 639.365 55.495 639.645 55.775 ;
        RECT 637.945 54.835 638.225 55.115 ;
        RECT 639.365 54.835 639.645 55.115 ;
        RECT 637.945 54.175 638.225 54.455 ;
        RECT 639.365 54.175 639.645 54.455 ;
        RECT 637.945 53.515 638.225 53.795 ;
        RECT 639.365 53.515 639.645 53.795 ;
        RECT 637.945 52.855 638.225 53.135 ;
        RECT 639.365 52.855 639.645 53.135 ;
        RECT 637.945 52.195 638.225 52.475 ;
        RECT 639.365 52.195 639.645 52.475 ;
        RECT 637.945 51.535 638.225 51.815 ;
        RECT 639.365 51.535 639.645 51.815 ;
        RECT 637.945 50.875 638.225 51.155 ;
        RECT 639.365 50.875 639.645 51.155 ;
        RECT 637.945 50.215 638.225 50.495 ;
        RECT 639.365 50.215 639.645 50.495 ;
        RECT 643.850 47.855 644.130 48.135 ;
        RECT 644.510 47.855 644.790 48.135 ;
        RECT 645.170 47.855 645.450 48.135 ;
        RECT 643.850 47.195 644.130 47.475 ;
        RECT 644.510 47.195 644.790 47.475 ;
        RECT 645.170 47.195 645.450 47.475 ;
        RECT 643.850 46.535 644.130 46.815 ;
        RECT 644.510 46.535 644.790 46.815 ;
        RECT 645.170 46.535 645.450 46.815 ;
        RECT 632.155 39.755 632.435 40.035 ;
        RECT 632.815 39.755 633.095 40.035 ;
        RECT 633.475 39.755 633.755 40.035 ;
        RECT 632.155 39.095 632.435 39.375 ;
        RECT 632.815 39.095 633.095 39.375 ;
        RECT 633.475 39.095 633.755 39.375 ;
        RECT 632.155 38.435 632.435 38.715 ;
        RECT 632.815 38.435 633.095 38.715 ;
        RECT 633.475 38.435 633.755 38.715 ;
        RECT 632.155 30.355 632.435 30.635 ;
        RECT 632.815 30.355 633.095 30.635 ;
        RECT 633.475 30.355 633.755 30.635 ;
        RECT 632.155 29.695 632.435 29.975 ;
        RECT 632.815 29.695 633.095 29.975 ;
        RECT 633.475 29.695 633.755 29.975 ;
        RECT 632.155 29.035 632.435 29.315 ;
        RECT 632.815 29.035 633.095 29.315 ;
        RECT 633.475 29.035 633.755 29.315 ;
        RECT 643.850 22.255 644.130 22.535 ;
        RECT 644.510 22.255 644.790 22.535 ;
        RECT 645.170 22.255 645.450 22.535 ;
        RECT 643.850 21.595 644.130 21.875 ;
        RECT 644.510 21.595 644.790 21.875 ;
        RECT 645.170 21.595 645.450 21.875 ;
        RECT 643.850 20.935 644.130 21.215 ;
        RECT 644.510 20.935 644.790 21.215 ;
        RECT 645.170 20.935 645.450 21.215 ;
        RECT 569.800 4.740 570.080 5.020 ;
        RECT 570.800 4.740 571.080 5.020 ;
        RECT 571.460 4.740 571.740 5.020 ;
        RECT 572.120 4.740 572.400 5.020 ;
        RECT 573.040 4.740 573.320 5.020 ;
        RECT 573.700 4.740 573.980 5.020 ;
        RECT 574.360 4.740 574.640 5.020 ;
        RECT 575.280 4.740 575.560 5.020 ;
        RECT 575.940 4.740 576.220 5.020 ;
        RECT 576.600 4.740 576.880 5.020 ;
        RECT 577.520 4.740 577.800 5.020 ;
        RECT 578.180 4.740 578.460 5.020 ;
        RECT 578.840 4.740 579.120 5.020 ;
        RECT 579.760 4.740 580.040 5.020 ;
        RECT 580.420 4.740 580.700 5.020 ;
        RECT 581.080 4.740 581.360 5.020 ;
        RECT 582.000 4.740 582.280 5.020 ;
        RECT 582.660 4.740 582.940 5.020 ;
        RECT 583.320 4.740 583.600 5.020 ;
        RECT 584.240 4.740 584.520 5.020 ;
        RECT 584.900 4.740 585.180 5.020 ;
        RECT 585.560 4.740 585.840 5.020 ;
        RECT 586.480 4.740 586.760 5.020 ;
        RECT 587.140 4.740 587.420 5.020 ;
        RECT 587.800 4.740 588.080 5.020 ;
        RECT 588.720 4.740 589.000 5.020 ;
        RECT 589.380 4.740 589.660 5.020 ;
        RECT 590.040 4.740 590.320 5.020 ;
        RECT 591.080 4.740 591.360 5.020 ;
        RECT 592.080 4.740 592.360 5.020 ;
        RECT 592.740 4.740 593.020 5.020 ;
        RECT 593.400 4.740 593.680 5.020 ;
        RECT 594.320 4.740 594.600 5.020 ;
        RECT 594.980 4.740 595.260 5.020 ;
        RECT 595.640 4.740 595.920 5.020 ;
        RECT 596.560 4.740 596.840 5.020 ;
        RECT 597.220 4.740 597.500 5.020 ;
        RECT 597.880 4.740 598.160 5.020 ;
        RECT 598.800 4.740 599.080 5.020 ;
        RECT 599.460 4.740 599.740 5.020 ;
        RECT 600.120 4.740 600.400 5.020 ;
        RECT 601.040 4.740 601.320 5.020 ;
        RECT 601.700 4.740 601.980 5.020 ;
        RECT 602.360 4.740 602.640 5.020 ;
        RECT 603.280 4.740 603.560 5.020 ;
        RECT 603.940 4.740 604.220 5.020 ;
        RECT 604.600 4.740 604.880 5.020 ;
        RECT 605.520 4.740 605.800 5.020 ;
        RECT 606.180 4.740 606.460 5.020 ;
        RECT 606.840 4.740 607.120 5.020 ;
        RECT 607.860 4.740 608.140 5.020 ;
        RECT 608.520 4.740 608.800 5.020 ;
        RECT 609.180 4.740 609.460 5.020 ;
        RECT 649.655 58.795 649.935 59.075 ;
        RECT 649.655 58.135 649.935 58.415 ;
        RECT 649.655 57.475 649.935 57.755 ;
        RECT 649.655 56.815 649.935 57.095 ;
        RECT 649.655 56.155 649.935 56.435 ;
        RECT 649.655 55.495 649.935 55.775 ;
        RECT 649.655 54.835 649.935 55.115 ;
        RECT 649.655 54.175 649.935 54.455 ;
        RECT 649.655 53.515 649.935 53.795 ;
        RECT 649.655 52.855 649.935 53.135 ;
        RECT 649.655 52.195 649.935 52.475 ;
        RECT 649.655 51.535 649.935 51.815 ;
        RECT 649.655 50.875 649.935 51.155 ;
        RECT 649.655 50.215 649.935 50.495 ;
        RECT 659.940 58.795 660.220 59.075 ;
        RECT 659.940 58.135 660.220 58.415 ;
        RECT 659.940 57.475 660.220 57.755 ;
        RECT 659.940 56.815 660.220 57.095 ;
        RECT 659.940 56.155 660.220 56.435 ;
        RECT 659.940 55.495 660.220 55.775 ;
        RECT 659.940 54.835 660.220 55.115 ;
        RECT 659.940 54.175 660.220 54.455 ;
        RECT 659.940 53.515 660.220 53.795 ;
        RECT 659.940 52.855 660.220 53.135 ;
        RECT 659.940 52.195 660.220 52.475 ;
        RECT 659.940 51.535 660.220 51.815 ;
        RECT 659.940 50.875 660.220 51.155 ;
        RECT 659.940 50.215 660.220 50.495 ;
        RECT 654.150 45.155 654.430 45.435 ;
        RECT 654.810 45.155 655.090 45.435 ;
        RECT 655.470 45.155 655.750 45.435 ;
        RECT 654.150 44.495 654.430 44.775 ;
        RECT 654.810 44.495 655.090 44.775 ;
        RECT 655.470 44.495 655.750 44.775 ;
        RECT 654.150 43.835 654.430 44.115 ;
        RECT 654.810 43.835 655.090 44.115 ;
        RECT 655.470 43.835 655.750 44.115 ;
        RECT 664.425 42.455 664.705 42.735 ;
        RECT 665.085 42.455 665.365 42.735 ;
        RECT 665.745 42.455 666.025 42.735 ;
        RECT 664.425 41.795 664.705 42.075 ;
        RECT 665.085 41.795 665.365 42.075 ;
        RECT 665.745 41.795 666.025 42.075 ;
        RECT 664.425 41.135 664.705 41.415 ;
        RECT 665.085 41.135 665.365 41.415 ;
        RECT 665.745 41.135 666.025 41.415 ;
        RECT 664.425 27.655 664.705 27.935 ;
        RECT 665.085 27.655 665.365 27.935 ;
        RECT 665.745 27.655 666.025 27.935 ;
        RECT 664.425 26.995 664.705 27.275 ;
        RECT 665.085 26.995 665.365 27.275 ;
        RECT 665.745 26.995 666.025 27.275 ;
        RECT 664.425 26.335 664.705 26.615 ;
        RECT 665.085 26.335 665.365 26.615 ;
        RECT 665.745 26.335 666.025 26.615 ;
        RECT 654.150 24.955 654.430 25.235 ;
        RECT 654.810 24.955 655.090 25.235 ;
        RECT 655.470 24.955 655.750 25.235 ;
        RECT 654.150 24.295 654.430 24.575 ;
        RECT 654.810 24.295 655.090 24.575 ;
        RECT 655.470 24.295 655.750 24.575 ;
        RECT 654.150 23.635 654.430 23.915 ;
        RECT 654.810 23.635 655.090 23.915 ;
        RECT 655.470 23.635 655.750 23.915 ;
        RECT 670.230 58.795 670.510 59.075 ;
        RECT 670.230 58.135 670.510 58.415 ;
        RECT 670.230 57.475 670.510 57.755 ;
        RECT 670.230 56.815 670.510 57.095 ;
        RECT 670.230 56.155 670.510 56.435 ;
        RECT 670.230 55.495 670.510 55.775 ;
        RECT 670.230 54.835 670.510 55.115 ;
        RECT 670.230 54.175 670.510 54.455 ;
        RECT 670.230 53.515 670.510 53.795 ;
        RECT 670.230 52.855 670.510 53.135 ;
        RECT 670.230 52.195 670.510 52.475 ;
        RECT 670.230 51.535 670.510 51.815 ;
        RECT 670.230 50.875 670.510 51.155 ;
        RECT 670.230 50.215 670.510 50.495 ;
        RECT 680.515 58.795 680.795 59.075 ;
        RECT 680.515 58.135 680.795 58.415 ;
        RECT 680.515 57.475 680.795 57.755 ;
        RECT 680.515 56.815 680.795 57.095 ;
        RECT 680.515 56.155 680.795 56.435 ;
        RECT 680.515 55.495 680.795 55.775 ;
        RECT 682.360 55.165 682.640 55.445 ;
        RECT 684.145 55.165 684.425 55.445 ;
        RECT 687.000 55.165 687.280 55.445 ;
        RECT 688.785 55.165 689.065 55.445 ;
        RECT 691.640 55.165 691.920 55.445 ;
        RECT 693.425 55.165 693.705 55.445 ;
        RECT 696.280 55.165 696.560 55.445 ;
        RECT 698.065 55.165 698.345 55.445 ;
        RECT 700.920 55.165 701.200 55.445 ;
        RECT 702.705 55.165 702.985 55.445 ;
        RECT 705.560 55.165 705.840 55.445 ;
        RECT 707.345 55.165 707.625 55.445 ;
        RECT 710.200 55.165 710.480 55.445 ;
        RECT 711.985 55.165 712.265 55.445 ;
        RECT 714.840 55.165 715.120 55.445 ;
        RECT 716.625 55.165 716.905 55.445 ;
        RECT 680.515 54.835 680.795 55.115 ;
        RECT 682.360 54.505 682.640 54.785 ;
        RECT 684.145 54.505 684.425 54.785 ;
        RECT 687.000 54.505 687.280 54.785 ;
        RECT 688.785 54.505 689.065 54.785 ;
        RECT 691.640 54.505 691.920 54.785 ;
        RECT 693.425 54.505 693.705 54.785 ;
        RECT 696.280 54.505 696.560 54.785 ;
        RECT 698.065 54.505 698.345 54.785 ;
        RECT 700.920 54.505 701.200 54.785 ;
        RECT 702.705 54.505 702.985 54.785 ;
        RECT 705.560 54.505 705.840 54.785 ;
        RECT 707.345 54.505 707.625 54.785 ;
        RECT 710.200 54.505 710.480 54.785 ;
        RECT 711.985 54.505 712.265 54.785 ;
        RECT 714.840 54.505 715.120 54.785 ;
        RECT 716.625 54.505 716.905 54.785 ;
        RECT 680.515 54.175 680.795 54.455 ;
        RECT 682.360 53.845 682.640 54.125 ;
        RECT 684.145 53.845 684.425 54.125 ;
        RECT 687.000 53.845 687.280 54.125 ;
        RECT 688.785 53.845 689.065 54.125 ;
        RECT 691.640 53.845 691.920 54.125 ;
        RECT 693.425 53.845 693.705 54.125 ;
        RECT 696.280 53.845 696.560 54.125 ;
        RECT 698.065 53.845 698.345 54.125 ;
        RECT 700.920 53.845 701.200 54.125 ;
        RECT 702.705 53.845 702.985 54.125 ;
        RECT 705.560 53.845 705.840 54.125 ;
        RECT 707.345 53.845 707.625 54.125 ;
        RECT 710.200 53.845 710.480 54.125 ;
        RECT 711.985 53.845 712.265 54.125 ;
        RECT 714.840 53.845 715.120 54.125 ;
        RECT 716.625 53.845 716.905 54.125 ;
        RECT 680.515 53.515 680.795 53.795 ;
        RECT 682.360 53.185 682.640 53.465 ;
        RECT 684.145 53.185 684.425 53.465 ;
        RECT 687.000 53.185 687.280 53.465 ;
        RECT 688.785 53.185 689.065 53.465 ;
        RECT 691.640 53.185 691.920 53.465 ;
        RECT 693.425 53.185 693.705 53.465 ;
        RECT 696.280 53.185 696.560 53.465 ;
        RECT 698.065 53.185 698.345 53.465 ;
        RECT 700.920 53.185 701.200 53.465 ;
        RECT 702.705 53.185 702.985 53.465 ;
        RECT 705.560 53.185 705.840 53.465 ;
        RECT 707.345 53.185 707.625 53.465 ;
        RECT 710.200 53.185 710.480 53.465 ;
        RECT 711.985 53.185 712.265 53.465 ;
        RECT 714.840 53.185 715.120 53.465 ;
        RECT 716.625 53.185 716.905 53.465 ;
        RECT 680.515 52.855 680.795 53.135 ;
        RECT 682.360 52.525 682.640 52.805 ;
        RECT 684.145 52.525 684.425 52.805 ;
        RECT 687.000 52.525 687.280 52.805 ;
        RECT 688.785 52.525 689.065 52.805 ;
        RECT 691.640 52.525 691.920 52.805 ;
        RECT 693.425 52.525 693.705 52.805 ;
        RECT 696.280 52.525 696.560 52.805 ;
        RECT 698.065 52.525 698.345 52.805 ;
        RECT 700.920 52.525 701.200 52.805 ;
        RECT 702.705 52.525 702.985 52.805 ;
        RECT 705.560 52.525 705.840 52.805 ;
        RECT 707.345 52.525 707.625 52.805 ;
        RECT 710.200 52.525 710.480 52.805 ;
        RECT 711.985 52.525 712.265 52.805 ;
        RECT 714.840 52.525 715.120 52.805 ;
        RECT 716.625 52.525 716.905 52.805 ;
        RECT 680.515 52.195 680.795 52.475 ;
        RECT 682.360 51.865 682.640 52.145 ;
        RECT 684.145 51.865 684.425 52.145 ;
        RECT 687.000 51.865 687.280 52.145 ;
        RECT 688.785 51.865 689.065 52.145 ;
        RECT 691.640 51.865 691.920 52.145 ;
        RECT 693.425 51.865 693.705 52.145 ;
        RECT 696.280 51.865 696.560 52.145 ;
        RECT 698.065 51.865 698.345 52.145 ;
        RECT 700.920 51.865 701.200 52.145 ;
        RECT 702.705 51.865 702.985 52.145 ;
        RECT 705.560 51.865 705.840 52.145 ;
        RECT 707.345 51.865 707.625 52.145 ;
        RECT 710.200 51.865 710.480 52.145 ;
        RECT 711.985 51.865 712.265 52.145 ;
        RECT 714.840 51.865 715.120 52.145 ;
        RECT 716.625 51.865 716.905 52.145 ;
        RECT 680.515 51.535 680.795 51.815 ;
        RECT 682.360 51.205 682.640 51.485 ;
        RECT 684.145 51.205 684.425 51.485 ;
        RECT 687.000 51.205 687.280 51.485 ;
        RECT 688.785 51.205 689.065 51.485 ;
        RECT 691.640 51.205 691.920 51.485 ;
        RECT 693.425 51.205 693.705 51.485 ;
        RECT 696.280 51.205 696.560 51.485 ;
        RECT 698.065 51.205 698.345 51.485 ;
        RECT 700.920 51.205 701.200 51.485 ;
        RECT 702.705 51.205 702.985 51.485 ;
        RECT 705.560 51.205 705.840 51.485 ;
        RECT 707.345 51.205 707.625 51.485 ;
        RECT 710.200 51.205 710.480 51.485 ;
        RECT 711.985 51.205 712.265 51.485 ;
        RECT 714.840 51.205 715.120 51.485 ;
        RECT 716.625 51.205 716.905 51.485 ;
        RECT 680.515 50.875 680.795 51.155 ;
        RECT 682.360 50.545 682.640 50.825 ;
        RECT 684.145 50.545 684.425 50.825 ;
        RECT 687.000 50.545 687.280 50.825 ;
        RECT 688.785 50.545 689.065 50.825 ;
        RECT 691.640 50.545 691.920 50.825 ;
        RECT 693.425 50.545 693.705 50.825 ;
        RECT 696.280 50.545 696.560 50.825 ;
        RECT 698.065 50.545 698.345 50.825 ;
        RECT 700.920 50.545 701.200 50.825 ;
        RECT 702.705 50.545 702.985 50.825 ;
        RECT 705.560 50.545 705.840 50.825 ;
        RECT 707.345 50.545 707.625 50.825 ;
        RECT 710.200 50.545 710.480 50.825 ;
        RECT 711.985 50.545 712.265 50.825 ;
        RECT 714.840 50.545 715.120 50.825 ;
        RECT 716.625 50.545 716.905 50.825 ;
        RECT 680.515 50.215 680.795 50.495 ;
        RECT 683.120 47.855 683.400 48.135 ;
        RECT 683.120 47.195 683.400 47.475 ;
        RECT 683.120 46.535 683.400 46.815 ;
        RECT 697.040 45.155 697.320 45.435 ;
        RECT 697.040 44.495 697.320 44.775 ;
        RECT 697.040 43.835 697.320 44.115 ;
        RECT 701.680 42.455 701.960 42.735 ;
        RECT 701.680 41.795 701.960 42.075 ;
        RECT 701.680 41.135 701.960 41.415 ;
        RECT 674.725 39.755 675.005 40.035 ;
        RECT 675.385 39.755 675.665 40.035 ;
        RECT 676.045 39.755 676.325 40.035 ;
        RECT 715.600 39.755 715.880 40.035 ;
        RECT 674.725 39.095 675.005 39.375 ;
        RECT 675.385 39.095 675.665 39.375 ;
        RECT 676.045 39.095 676.325 39.375 ;
        RECT 715.600 39.095 715.880 39.375 ;
        RECT 674.725 38.435 675.005 38.715 ;
        RECT 675.385 38.435 675.665 38.715 ;
        RECT 676.045 38.435 676.325 38.715 ;
        RECT 715.600 38.435 715.880 38.715 ;
        RECT 674.725 30.355 675.005 30.635 ;
        RECT 675.385 30.355 675.665 30.635 ;
        RECT 676.045 30.355 676.325 30.635 ;
        RECT 710.960 30.355 711.240 30.635 ;
        RECT 674.725 29.695 675.005 29.975 ;
        RECT 675.385 29.695 675.665 29.975 ;
        RECT 676.045 29.695 676.325 29.975 ;
        RECT 710.960 29.695 711.240 29.975 ;
        RECT 674.725 29.035 675.005 29.315 ;
        RECT 675.385 29.035 675.665 29.315 ;
        RECT 676.045 29.035 676.325 29.315 ;
        RECT 710.960 29.035 711.240 29.315 ;
        RECT 706.320 27.655 706.600 27.935 ;
        RECT 706.320 26.995 706.600 27.275 ;
        RECT 706.320 26.335 706.600 26.615 ;
        RECT 692.400 24.955 692.680 25.235 ;
        RECT 692.400 24.295 692.680 24.575 ;
        RECT 692.400 23.635 692.680 23.915 ;
        RECT 687.760 22.255 688.040 22.535 ;
        RECT 687.760 21.595 688.040 21.875 ;
        RECT 687.760 20.935 688.040 21.215 ;
        RECT 682.360 18.165 682.640 18.445 ;
        RECT 684.145 18.165 684.425 18.445 ;
        RECT 687.000 18.165 687.280 18.445 ;
        RECT 688.785 18.165 689.065 18.445 ;
        RECT 691.640 18.165 691.920 18.445 ;
        RECT 693.425 18.165 693.705 18.445 ;
        RECT 696.280 18.165 696.560 18.445 ;
        RECT 698.065 18.165 698.345 18.445 ;
        RECT 700.920 18.165 701.200 18.445 ;
        RECT 702.705 18.165 702.985 18.445 ;
        RECT 705.560 18.165 705.840 18.445 ;
        RECT 707.345 18.165 707.625 18.445 ;
        RECT 710.200 18.165 710.480 18.445 ;
        RECT 711.985 18.165 712.265 18.445 ;
        RECT 714.840 18.165 715.120 18.445 ;
        RECT 716.625 18.165 716.905 18.445 ;
        RECT 682.360 17.505 682.640 17.785 ;
        RECT 684.145 17.505 684.425 17.785 ;
        RECT 687.000 17.505 687.280 17.785 ;
        RECT 688.785 17.505 689.065 17.785 ;
        RECT 691.640 17.505 691.920 17.785 ;
        RECT 693.425 17.505 693.705 17.785 ;
        RECT 696.280 17.505 696.560 17.785 ;
        RECT 698.065 17.505 698.345 17.785 ;
        RECT 700.920 17.505 701.200 17.785 ;
        RECT 702.705 17.505 702.985 17.785 ;
        RECT 705.560 17.505 705.840 17.785 ;
        RECT 707.345 17.505 707.625 17.785 ;
        RECT 710.200 17.505 710.480 17.785 ;
        RECT 711.985 17.505 712.265 17.785 ;
        RECT 714.840 17.505 715.120 17.785 ;
        RECT 716.625 17.505 716.905 17.785 ;
        RECT 682.360 16.845 682.640 17.125 ;
        RECT 684.145 16.845 684.425 17.125 ;
        RECT 687.000 16.845 687.280 17.125 ;
        RECT 688.785 16.845 689.065 17.125 ;
        RECT 691.640 16.845 691.920 17.125 ;
        RECT 693.425 16.845 693.705 17.125 ;
        RECT 696.280 16.845 696.560 17.125 ;
        RECT 698.065 16.845 698.345 17.125 ;
        RECT 700.920 16.845 701.200 17.125 ;
        RECT 702.705 16.845 702.985 17.125 ;
        RECT 705.560 16.845 705.840 17.125 ;
        RECT 707.345 16.845 707.625 17.125 ;
        RECT 710.200 16.845 710.480 17.125 ;
        RECT 711.985 16.845 712.265 17.125 ;
        RECT 714.840 16.845 715.120 17.125 ;
        RECT 716.625 16.845 716.905 17.125 ;
        RECT 682.360 16.185 682.640 16.465 ;
        RECT 684.145 16.185 684.425 16.465 ;
        RECT 687.000 16.185 687.280 16.465 ;
        RECT 688.785 16.185 689.065 16.465 ;
        RECT 691.640 16.185 691.920 16.465 ;
        RECT 693.425 16.185 693.705 16.465 ;
        RECT 696.280 16.185 696.560 16.465 ;
        RECT 698.065 16.185 698.345 16.465 ;
        RECT 700.920 16.185 701.200 16.465 ;
        RECT 702.705 16.185 702.985 16.465 ;
        RECT 705.560 16.185 705.840 16.465 ;
        RECT 707.345 16.185 707.625 16.465 ;
        RECT 710.200 16.185 710.480 16.465 ;
        RECT 711.985 16.185 712.265 16.465 ;
        RECT 714.840 16.185 715.120 16.465 ;
        RECT 716.625 16.185 716.905 16.465 ;
        RECT 682.360 15.525 682.640 15.805 ;
        RECT 684.145 15.525 684.425 15.805 ;
        RECT 687.000 15.525 687.280 15.805 ;
        RECT 688.785 15.525 689.065 15.805 ;
        RECT 691.640 15.525 691.920 15.805 ;
        RECT 693.425 15.525 693.705 15.805 ;
        RECT 696.280 15.525 696.560 15.805 ;
        RECT 698.065 15.525 698.345 15.805 ;
        RECT 700.920 15.525 701.200 15.805 ;
        RECT 702.705 15.525 702.985 15.805 ;
        RECT 705.560 15.525 705.840 15.805 ;
        RECT 707.345 15.525 707.625 15.805 ;
        RECT 710.200 15.525 710.480 15.805 ;
        RECT 711.985 15.525 712.265 15.805 ;
        RECT 714.840 15.525 715.120 15.805 ;
        RECT 716.625 15.525 716.905 15.805 ;
        RECT 682.360 14.865 682.640 15.145 ;
        RECT 684.145 14.865 684.425 15.145 ;
        RECT 687.000 14.865 687.280 15.145 ;
        RECT 688.785 14.865 689.065 15.145 ;
        RECT 691.640 14.865 691.920 15.145 ;
        RECT 693.425 14.865 693.705 15.145 ;
        RECT 696.280 14.865 696.560 15.145 ;
        RECT 698.065 14.865 698.345 15.145 ;
        RECT 700.920 14.865 701.200 15.145 ;
        RECT 702.705 14.865 702.985 15.145 ;
        RECT 705.560 14.865 705.840 15.145 ;
        RECT 707.345 14.865 707.625 15.145 ;
        RECT 710.200 14.865 710.480 15.145 ;
        RECT 711.985 14.865 712.265 15.145 ;
        RECT 714.840 14.865 715.120 15.145 ;
        RECT 716.625 14.865 716.905 15.145 ;
        RECT 682.360 14.205 682.640 14.485 ;
        RECT 684.145 14.205 684.425 14.485 ;
        RECT 687.000 14.205 687.280 14.485 ;
        RECT 688.785 14.205 689.065 14.485 ;
        RECT 691.640 14.205 691.920 14.485 ;
        RECT 693.425 14.205 693.705 14.485 ;
        RECT 696.280 14.205 696.560 14.485 ;
        RECT 698.065 14.205 698.345 14.485 ;
        RECT 700.920 14.205 701.200 14.485 ;
        RECT 702.705 14.205 702.985 14.485 ;
        RECT 705.560 14.205 705.840 14.485 ;
        RECT 707.345 14.205 707.625 14.485 ;
        RECT 710.200 14.205 710.480 14.485 ;
        RECT 711.985 14.205 712.265 14.485 ;
        RECT 714.840 14.205 715.120 14.485 ;
        RECT 716.625 14.205 716.905 14.485 ;
        RECT 682.360 13.545 682.640 13.825 ;
        RECT 684.145 13.545 684.425 13.825 ;
        RECT 687.000 13.545 687.280 13.825 ;
        RECT 688.785 13.545 689.065 13.825 ;
        RECT 691.640 13.545 691.920 13.825 ;
        RECT 693.425 13.545 693.705 13.825 ;
        RECT 696.280 13.545 696.560 13.825 ;
        RECT 698.065 13.545 698.345 13.825 ;
        RECT 700.920 13.545 701.200 13.825 ;
        RECT 702.705 13.545 702.985 13.825 ;
        RECT 705.560 13.545 705.840 13.825 ;
        RECT 707.345 13.545 707.625 13.825 ;
        RECT 710.200 13.545 710.480 13.825 ;
        RECT 711.985 13.545 712.265 13.825 ;
        RECT 714.840 13.545 715.120 13.825 ;
        RECT 716.625 13.545 716.905 13.825 ;
        RECT 682.360 12.885 682.640 13.165 ;
        RECT 684.145 12.885 684.425 13.165 ;
        RECT 687.000 12.885 687.280 13.165 ;
        RECT 688.785 12.885 689.065 13.165 ;
        RECT 691.640 12.885 691.920 13.165 ;
        RECT 693.425 12.885 693.705 13.165 ;
        RECT 696.280 12.885 696.560 13.165 ;
        RECT 698.065 12.885 698.345 13.165 ;
        RECT 700.920 12.885 701.200 13.165 ;
        RECT 702.705 12.885 702.985 13.165 ;
        RECT 705.560 12.885 705.840 13.165 ;
        RECT 707.345 12.885 707.625 13.165 ;
        RECT 710.200 12.885 710.480 13.165 ;
        RECT 711.985 12.885 712.265 13.165 ;
        RECT 714.840 12.885 715.120 13.165 ;
        RECT 716.625 12.885 716.905 13.165 ;
        RECT 682.360 12.225 682.640 12.505 ;
        RECT 684.145 12.225 684.425 12.505 ;
        RECT 687.000 12.225 687.280 12.505 ;
        RECT 688.785 12.225 689.065 12.505 ;
        RECT 691.640 12.225 691.920 12.505 ;
        RECT 693.425 12.225 693.705 12.505 ;
        RECT 696.280 12.225 696.560 12.505 ;
        RECT 698.065 12.225 698.345 12.505 ;
        RECT 700.920 12.225 701.200 12.505 ;
        RECT 702.705 12.225 702.985 12.505 ;
        RECT 705.560 12.225 705.840 12.505 ;
        RECT 707.345 12.225 707.625 12.505 ;
        RECT 710.200 12.225 710.480 12.505 ;
        RECT 711.985 12.225 712.265 12.505 ;
        RECT 714.840 12.225 715.120 12.505 ;
        RECT 716.625 12.225 716.905 12.505 ;
        RECT 682.360 11.565 682.640 11.845 ;
        RECT 684.145 11.565 684.425 11.845 ;
        RECT 687.000 11.565 687.280 11.845 ;
        RECT 688.785 11.565 689.065 11.845 ;
        RECT 691.640 11.565 691.920 11.845 ;
        RECT 693.425 11.565 693.705 11.845 ;
        RECT 696.280 11.565 696.560 11.845 ;
        RECT 698.065 11.565 698.345 11.845 ;
        RECT 700.920 11.565 701.200 11.845 ;
        RECT 702.705 11.565 702.985 11.845 ;
        RECT 705.560 11.565 705.840 11.845 ;
        RECT 707.345 11.565 707.625 11.845 ;
        RECT 710.200 11.565 710.480 11.845 ;
        RECT 711.985 11.565 712.265 11.845 ;
        RECT 714.840 11.565 715.120 11.845 ;
        RECT 716.625 11.565 716.905 11.845 ;
        RECT 682.360 10.905 682.640 11.185 ;
        RECT 684.145 10.905 684.425 11.185 ;
        RECT 687.000 10.905 687.280 11.185 ;
        RECT 688.785 10.905 689.065 11.185 ;
        RECT 691.640 10.905 691.920 11.185 ;
        RECT 693.425 10.905 693.705 11.185 ;
        RECT 696.280 10.905 696.560 11.185 ;
        RECT 698.065 10.905 698.345 11.185 ;
        RECT 700.920 10.905 701.200 11.185 ;
        RECT 702.705 10.905 702.985 11.185 ;
        RECT 705.560 10.905 705.840 11.185 ;
        RECT 707.345 10.905 707.625 11.185 ;
        RECT 710.200 10.905 710.480 11.185 ;
        RECT 711.985 10.905 712.265 11.185 ;
        RECT 714.840 10.905 715.120 11.185 ;
        RECT 716.625 10.905 716.905 11.185 ;
        RECT 682.360 10.245 682.640 10.525 ;
        RECT 684.145 10.245 684.425 10.525 ;
        RECT 687.000 10.245 687.280 10.525 ;
        RECT 688.785 10.245 689.065 10.525 ;
        RECT 691.640 10.245 691.920 10.525 ;
        RECT 693.425 10.245 693.705 10.525 ;
        RECT 696.280 10.245 696.560 10.525 ;
        RECT 698.065 10.245 698.345 10.525 ;
        RECT 700.920 10.245 701.200 10.525 ;
        RECT 702.705 10.245 702.985 10.525 ;
        RECT 705.560 10.245 705.840 10.525 ;
        RECT 707.345 10.245 707.625 10.525 ;
        RECT 710.200 10.245 710.480 10.525 ;
        RECT 711.985 10.245 712.265 10.525 ;
        RECT 714.840 10.245 715.120 10.525 ;
        RECT 716.625 10.245 716.905 10.525 ;
        RECT 682.360 9.585 682.640 9.865 ;
        RECT 684.145 9.585 684.425 9.865 ;
        RECT 687.000 9.585 687.280 9.865 ;
        RECT 688.785 9.585 689.065 9.865 ;
        RECT 691.640 9.585 691.920 9.865 ;
        RECT 693.425 9.585 693.705 9.865 ;
        RECT 696.280 9.585 696.560 9.865 ;
        RECT 698.065 9.585 698.345 9.865 ;
        RECT 700.920 9.585 701.200 9.865 ;
        RECT 702.705 9.585 702.985 9.865 ;
        RECT 705.560 9.585 705.840 9.865 ;
        RECT 707.345 9.585 707.625 9.865 ;
        RECT 710.200 9.585 710.480 9.865 ;
        RECT 711.985 9.585 712.265 9.865 ;
        RECT 714.840 9.585 715.120 9.865 ;
        RECT 716.625 9.585 716.905 9.865 ;
        RECT 611.240 4.740 611.520 5.020 ;
        RECT 612.240 4.740 612.520 5.020 ;
        RECT 612.900 4.740 613.180 5.020 ;
        RECT 613.560 4.740 613.840 5.020 ;
        RECT 614.480 4.740 614.760 5.020 ;
        RECT 615.140 4.740 615.420 5.020 ;
        RECT 615.800 4.740 616.080 5.020 ;
        RECT 616.720 4.740 617.000 5.020 ;
        RECT 617.380 4.740 617.660 5.020 ;
        RECT 618.040 4.740 618.320 5.020 ;
        RECT 618.960 4.740 619.240 5.020 ;
        RECT 619.620 4.740 619.900 5.020 ;
        RECT 620.280 4.740 620.560 5.020 ;
        RECT 621.200 4.740 621.480 5.020 ;
        RECT 621.860 4.740 622.140 5.020 ;
        RECT 622.520 4.740 622.800 5.020 ;
        RECT 623.440 4.740 623.720 5.020 ;
        RECT 624.100 4.740 624.380 5.020 ;
        RECT 624.760 4.740 625.040 5.020 ;
        RECT 625.680 4.740 625.960 5.020 ;
        RECT 626.340 4.740 626.620 5.020 ;
        RECT 627.000 4.740 627.280 5.020 ;
        RECT 627.920 4.740 628.200 5.020 ;
        RECT 628.580 4.740 628.860 5.020 ;
        RECT 629.240 4.740 629.520 5.020 ;
        RECT 630.160 4.740 630.440 5.020 ;
        RECT 630.820 4.740 631.100 5.020 ;
        RECT 631.480 4.740 631.760 5.020 ;
        RECT 632.520 4.740 632.800 5.020 ;
        RECT 633.520 4.740 633.800 5.020 ;
        RECT 634.180 4.740 634.460 5.020 ;
        RECT 634.840 4.740 635.120 5.020 ;
        RECT 635.760 4.740 636.040 5.020 ;
        RECT 636.420 4.740 636.700 5.020 ;
        RECT 637.080 4.740 637.360 5.020 ;
        RECT 638.000 4.740 638.280 5.020 ;
        RECT 638.660 4.740 638.940 5.020 ;
        RECT 639.320 4.740 639.600 5.020 ;
        RECT 640.240 4.740 640.520 5.020 ;
        RECT 640.900 4.740 641.180 5.020 ;
        RECT 641.560 4.740 641.840 5.020 ;
        RECT 642.480 4.740 642.760 5.020 ;
        RECT 643.140 4.740 643.420 5.020 ;
        RECT 643.800 4.740 644.080 5.020 ;
        RECT 644.720 4.740 645.000 5.020 ;
        RECT 645.380 4.740 645.660 5.020 ;
        RECT 646.040 4.740 646.320 5.020 ;
        RECT 646.960 4.740 647.240 5.020 ;
        RECT 647.620 4.740 647.900 5.020 ;
        RECT 648.280 4.740 648.560 5.020 ;
        RECT 649.200 4.740 649.480 5.020 ;
        RECT 649.860 4.740 650.140 5.020 ;
        RECT 650.520 4.740 650.800 5.020 ;
        RECT 651.540 4.740 651.820 5.020 ;
        RECT 652.200 4.740 652.480 5.020 ;
        RECT 652.860 4.740 653.140 5.020 ;
        RECT 682.360 8.925 682.640 9.205 ;
        RECT 684.145 8.925 684.425 9.205 ;
        RECT 687.000 8.925 687.280 9.205 ;
        RECT 688.785 8.925 689.065 9.205 ;
        RECT 691.640 8.925 691.920 9.205 ;
        RECT 693.425 8.925 693.705 9.205 ;
        RECT 696.280 8.925 696.560 9.205 ;
        RECT 698.065 8.925 698.345 9.205 ;
        RECT 700.920 8.925 701.200 9.205 ;
        RECT 702.705 8.925 702.985 9.205 ;
        RECT 705.560 8.925 705.840 9.205 ;
        RECT 707.345 8.925 707.625 9.205 ;
        RECT 710.200 8.925 710.480 9.205 ;
        RECT 711.985 8.925 712.265 9.205 ;
        RECT 714.840 8.925 715.120 9.205 ;
        RECT 716.625 8.925 716.905 9.205 ;
        RECT 654.920 4.740 655.200 5.020 ;
        RECT 655.920 4.740 656.200 5.020 ;
        RECT 656.580 4.740 656.860 5.020 ;
        RECT 657.240 4.740 657.520 5.020 ;
        RECT 658.160 4.740 658.440 5.020 ;
        RECT 658.820 4.740 659.100 5.020 ;
        RECT 659.480 4.740 659.760 5.020 ;
        RECT 660.400 4.740 660.680 5.020 ;
        RECT 661.060 4.740 661.340 5.020 ;
        RECT 661.720 4.740 662.000 5.020 ;
        RECT 662.640 4.740 662.920 5.020 ;
        RECT 663.300 4.740 663.580 5.020 ;
        RECT 663.960 4.740 664.240 5.020 ;
        RECT 664.880 4.740 665.160 5.020 ;
        RECT 665.540 4.740 665.820 5.020 ;
        RECT 666.200 4.740 666.480 5.020 ;
        RECT 667.120 4.740 667.400 5.020 ;
        RECT 667.780 4.740 668.060 5.020 ;
        RECT 668.440 4.740 668.720 5.020 ;
        RECT 669.360 4.740 669.640 5.020 ;
        RECT 670.020 4.740 670.300 5.020 ;
        RECT 670.680 4.740 670.960 5.020 ;
        RECT 671.600 4.740 671.880 5.020 ;
        RECT 672.260 4.740 672.540 5.020 ;
        RECT 672.920 4.740 673.200 5.020 ;
        RECT 673.840 4.740 674.120 5.020 ;
        RECT 674.500 4.740 674.780 5.020 ;
        RECT 675.160 4.740 675.440 5.020 ;
        RECT 676.200 4.740 676.480 5.020 ;
        RECT 677.200 4.740 677.480 5.020 ;
        RECT 677.860 4.740 678.140 5.020 ;
        RECT 678.520 4.740 678.800 5.020 ;
        RECT 679.540 4.740 679.820 5.020 ;
        RECT 121.470 3.470 121.750 3.750 ;
        RECT 121.880 2.810 122.160 3.090 ;
        RECT 0.900 0.820 1.180 1.100 ;
        RECT 2.040 0.820 2.320 1.100 ;
        RECT 7.480 0.820 7.760 1.100 ;
        RECT 8.140 0.820 8.420 1.100 ;
        RECT 8.800 0.820 9.080 1.100 ;
        RECT 14.350 0.820 14.630 1.100 ;
        RECT 15.670 0.820 15.950 1.100 ;
        RECT 17.710 0.820 17.990 1.100 ;
        RECT 19.030 0.820 19.310 1.100 ;
        RECT 25.670 0.820 25.950 1.100 ;
        RECT 26.330 0.820 26.610 1.100 ;
        RECT 26.990 0.820 27.270 1.100 ;
        RECT 32.540 0.820 32.820 1.100 ;
        RECT 33.860 0.820 34.140 1.100 ;
        RECT 36.180 0.820 36.460 1.100 ;
        RECT 41.620 0.820 41.900 1.100 ;
        RECT 42.280 0.820 42.560 1.100 ;
        RECT 42.940 0.820 43.220 1.100 ;
        RECT 48.490 0.820 48.770 1.100 ;
        RECT 49.810 0.820 50.090 1.100 ;
        RECT 56.450 0.820 56.730 1.100 ;
        RECT 57.110 0.820 57.390 1.100 ;
        RECT 57.770 0.820 58.050 1.100 ;
        RECT 63.320 0.820 63.600 1.100 ;
        RECT 64.640 0.820 64.920 1.100 ;
        RECT 66.680 0.820 66.960 1.100 ;
        RECT 68.000 0.820 68.280 1.100 ;
        RECT 70.320 0.820 70.600 1.100 ;
        RECT 75.760 0.820 76.040 1.100 ;
        RECT 76.420 0.820 76.700 1.100 ;
        RECT 77.080 0.820 77.360 1.100 ;
        RECT 82.630 0.820 82.910 1.100 ;
        RECT 83.950 0.820 84.230 1.100 ;
        RECT 90.590 0.820 90.870 1.100 ;
        RECT 91.250 0.820 91.530 1.100 ;
        RECT 91.910 0.820 92.190 1.100 ;
        RECT 97.460 0.820 97.740 1.100 ;
        RECT 98.780 0.820 99.060 1.100 ;
        RECT 100.820 0.820 101.100 1.100 ;
        RECT 102.140 0.820 102.420 1.100 ;
        RECT 104.460 0.820 104.740 1.100 ;
        RECT 109.900 0.820 110.180 1.100 ;
        RECT 110.560 0.820 110.840 1.100 ;
        RECT 111.220 0.820 111.500 1.100 ;
        RECT 116.770 0.820 117.050 1.100 ;
        RECT 118.090 0.820 118.370 1.100 ;
        RECT 124.730 0.820 125.010 1.100 ;
        RECT 125.390 0.820 125.670 1.100 ;
        RECT 126.050 0.820 126.330 1.100 ;
        RECT 131.600 0.820 131.880 1.100 ;
        RECT 132.920 0.820 133.200 1.100 ;
        RECT 135.240 0.820 135.520 1.100 ;
        RECT 136.240 0.820 136.520 1.100 ;
        RECT 136.900 0.820 137.180 1.100 ;
        RECT 137.560 0.820 137.840 1.100 ;
        RECT 138.480 0.820 138.760 1.100 ;
        RECT 139.140 0.820 139.420 1.100 ;
        RECT 139.800 0.820 140.080 1.100 ;
        RECT 140.560 0.820 140.840 1.100 ;
        RECT 141.880 0.820 142.160 1.100 ;
        RECT 144.080 0.820 144.360 1.100 ;
        RECT 144.740 0.820 145.020 1.100 ;
        RECT 145.400 0.820 145.680 1.100 ;
        RECT 146.320 0.820 146.600 1.100 ;
        RECT 146.980 0.820 147.260 1.100 ;
        RECT 147.640 0.820 147.920 1.100 ;
        RECT 148.560 0.820 148.840 1.100 ;
        RECT 149.220 0.820 149.500 1.100 ;
        RECT 149.880 0.820 150.160 1.100 ;
        RECT 150.800 0.820 151.080 1.100 ;
        RECT 151.460 0.820 151.740 1.100 ;
        RECT 152.120 0.820 152.400 1.100 ;
        RECT 153.040 0.820 153.320 1.100 ;
        RECT 153.700 0.820 153.980 1.100 ;
        RECT 154.360 0.820 154.640 1.100 ;
        RECT 155.400 0.820 155.680 1.100 ;
        RECT 156.400 0.820 156.680 1.100 ;
        RECT 157.060 0.820 157.340 1.100 ;
        RECT 157.720 0.820 158.000 1.100 ;
        RECT 158.640 0.820 158.920 1.100 ;
        RECT 159.300 0.820 159.580 1.100 ;
        RECT 159.960 0.820 160.240 1.100 ;
        RECT 160.880 0.820 161.160 1.100 ;
        RECT 161.540 0.820 161.820 1.100 ;
        RECT 162.200 0.820 162.480 1.100 ;
        RECT 163.120 0.820 163.400 1.100 ;
        RECT 163.780 0.820 164.060 1.100 ;
        RECT 164.440 0.820 164.720 1.100 ;
        RECT 165.360 0.820 165.640 1.100 ;
        RECT 166.020 0.820 166.300 1.100 ;
        RECT 166.680 0.820 166.960 1.100 ;
        RECT 167.600 0.820 167.880 1.100 ;
        RECT 168.260 0.820 168.540 1.100 ;
        RECT 168.920 0.820 169.200 1.100 ;
        RECT 169.840 0.820 170.120 1.100 ;
        RECT 170.500 0.820 170.780 1.100 ;
        RECT 171.160 0.820 171.440 1.100 ;
        RECT 172.080 0.820 172.360 1.100 ;
        RECT 172.740 0.820 173.020 1.100 ;
        RECT 173.400 0.820 173.680 1.100 ;
        RECT 174.320 0.820 174.600 1.100 ;
        RECT 174.980 0.820 175.260 1.100 ;
        RECT 175.640 0.820 175.920 1.100 ;
        RECT 176.680 0.820 176.960 1.100 ;
        RECT 177.680 0.820 177.960 1.100 ;
        RECT 178.340 0.820 178.620 1.100 ;
        RECT 179.000 0.820 179.280 1.100 ;
        RECT 179.920 0.820 180.200 1.100 ;
        RECT 180.580 0.820 180.860 1.100 ;
        RECT 181.240 0.820 181.520 1.100 ;
        RECT 182.000 0.820 182.280 1.100 ;
        RECT 183.320 0.820 183.600 1.100 ;
        RECT 185.520 0.820 185.800 1.100 ;
        RECT 186.180 0.820 186.460 1.100 ;
        RECT 186.840 0.820 187.120 1.100 ;
        RECT 187.760 0.820 188.040 1.100 ;
        RECT 188.420 0.820 188.700 1.100 ;
        RECT 189.080 0.820 189.360 1.100 ;
        RECT 190.000 0.820 190.280 1.100 ;
        RECT 190.660 0.820 190.940 1.100 ;
        RECT 191.320 0.820 191.600 1.100 ;
        RECT 192.240 0.820 192.520 1.100 ;
        RECT 192.900 0.820 193.180 1.100 ;
        RECT 193.560 0.820 193.840 1.100 ;
        RECT 194.480 0.820 194.760 1.100 ;
        RECT 195.140 0.820 195.420 1.100 ;
        RECT 195.800 0.820 196.080 1.100 ;
        RECT 196.840 0.820 197.120 1.100 ;
        RECT 197.840 0.820 198.120 1.100 ;
        RECT 198.500 0.820 198.780 1.100 ;
        RECT 199.160 0.820 199.440 1.100 ;
        RECT 200.080 0.820 200.360 1.100 ;
        RECT 200.740 0.820 201.020 1.100 ;
        RECT 201.400 0.820 201.680 1.100 ;
        RECT 202.320 0.820 202.600 1.100 ;
        RECT 202.980 0.820 203.260 1.100 ;
        RECT 203.640 0.820 203.920 1.100 ;
        RECT 204.560 0.820 204.840 1.100 ;
        RECT 205.220 0.820 205.500 1.100 ;
        RECT 205.880 0.820 206.160 1.100 ;
        RECT 206.800 0.820 207.080 1.100 ;
        RECT 207.460 0.820 207.740 1.100 ;
        RECT 208.120 0.820 208.400 1.100 ;
        RECT 209.040 0.820 209.320 1.100 ;
        RECT 209.700 0.820 209.980 1.100 ;
        RECT 210.360 0.820 210.640 1.100 ;
        RECT 211.280 0.820 211.560 1.100 ;
        RECT 211.940 0.820 212.220 1.100 ;
        RECT 212.600 0.820 212.880 1.100 ;
        RECT 213.520 0.820 213.800 1.100 ;
        RECT 214.180 0.820 214.460 1.100 ;
        RECT 214.840 0.820 215.120 1.100 ;
        RECT 215.760 0.820 216.040 1.100 ;
        RECT 216.420 0.820 216.700 1.100 ;
        RECT 217.080 0.820 217.360 1.100 ;
        RECT 218.120 0.820 218.400 1.100 ;
        RECT 219.120 0.820 219.400 1.100 ;
        RECT 219.780 0.820 220.060 1.100 ;
        RECT 220.440 0.820 220.720 1.100 ;
        RECT 221.360 0.820 221.640 1.100 ;
        RECT 222.020 0.820 222.300 1.100 ;
        RECT 222.680 0.820 222.960 1.100 ;
        RECT 223.600 0.820 223.880 1.100 ;
        RECT 224.260 0.820 224.540 1.100 ;
        RECT 224.920 0.820 225.200 1.100 ;
        RECT 225.680 0.820 225.960 1.100 ;
        RECT 227.000 0.820 227.280 1.100 ;
        RECT 229.200 0.820 229.480 1.100 ;
        RECT 229.860 0.820 230.140 1.100 ;
        RECT 230.520 0.820 230.800 1.100 ;
        RECT 231.440 0.820 231.720 1.100 ;
        RECT 232.100 0.820 232.380 1.100 ;
        RECT 232.760 0.820 233.040 1.100 ;
        RECT 233.680 0.820 233.960 1.100 ;
        RECT 234.340 0.820 234.620 1.100 ;
        RECT 235.000 0.820 235.280 1.100 ;
        RECT 235.920 0.820 236.200 1.100 ;
        RECT 236.580 0.820 236.860 1.100 ;
        RECT 237.240 0.820 237.520 1.100 ;
        RECT 238.280 0.820 238.560 1.100 ;
        RECT 239.280 0.820 239.560 1.100 ;
        RECT 239.940 0.820 240.220 1.100 ;
        RECT 240.600 0.820 240.880 1.100 ;
        RECT 241.520 0.820 241.800 1.100 ;
        RECT 242.180 0.820 242.460 1.100 ;
        RECT 242.840 0.820 243.120 1.100 ;
        RECT 243.760 0.820 244.040 1.100 ;
        RECT 244.420 0.820 244.700 1.100 ;
        RECT 245.080 0.820 245.360 1.100 ;
        RECT 246.000 0.820 246.280 1.100 ;
        RECT 246.660 0.820 246.940 1.100 ;
        RECT 247.320 0.820 247.600 1.100 ;
        RECT 248.240 0.820 248.520 1.100 ;
        RECT 248.900 0.820 249.180 1.100 ;
        RECT 249.560 0.820 249.840 1.100 ;
        RECT 250.480 0.820 250.760 1.100 ;
        RECT 251.140 0.820 251.420 1.100 ;
        RECT 251.800 0.820 252.080 1.100 ;
        RECT 252.720 0.820 253.000 1.100 ;
        RECT 253.380 0.820 253.660 1.100 ;
        RECT 254.040 0.820 254.320 1.100 ;
        RECT 254.960 0.820 255.240 1.100 ;
        RECT 255.620 0.820 255.900 1.100 ;
        RECT 256.280 0.820 256.560 1.100 ;
        RECT 257.200 0.820 257.480 1.100 ;
        RECT 257.860 0.820 258.140 1.100 ;
        RECT 258.520 0.820 258.800 1.100 ;
        RECT 259.560 0.820 259.840 1.100 ;
        RECT 260.560 0.820 260.840 1.100 ;
        RECT 261.220 0.820 261.500 1.100 ;
        RECT 261.880 0.820 262.160 1.100 ;
        RECT 262.800 0.820 263.080 1.100 ;
        RECT 263.460 0.820 263.740 1.100 ;
        RECT 264.120 0.820 264.400 1.100 ;
        RECT 265.040 0.820 265.320 1.100 ;
        RECT 265.700 0.820 265.980 1.100 ;
        RECT 266.360 0.820 266.640 1.100 ;
        RECT 267.120 0.820 267.400 1.100 ;
        RECT 268.440 0.820 268.720 1.100 ;
        RECT 270.640 0.820 270.920 1.100 ;
        RECT 271.300 0.820 271.580 1.100 ;
        RECT 271.960 0.820 272.240 1.100 ;
        RECT 272.880 0.820 273.160 1.100 ;
        RECT 273.540 0.820 273.820 1.100 ;
        RECT 274.200 0.820 274.480 1.100 ;
        RECT 275.120 0.820 275.400 1.100 ;
        RECT 275.780 0.820 276.060 1.100 ;
        RECT 276.440 0.820 276.720 1.100 ;
        RECT 277.360 0.820 277.640 1.100 ;
        RECT 278.020 0.820 278.300 1.100 ;
        RECT 278.680 0.820 278.960 1.100 ;
        RECT 279.720 0.820 280.000 1.100 ;
        RECT 280.720 0.820 281.000 1.100 ;
        RECT 281.380 0.820 281.660 1.100 ;
        RECT 282.040 0.820 282.320 1.100 ;
        RECT 282.960 0.820 283.240 1.100 ;
        RECT 283.620 0.820 283.900 1.100 ;
        RECT 284.280 0.820 284.560 1.100 ;
        RECT 285.200 0.820 285.480 1.100 ;
        RECT 285.860 0.820 286.140 1.100 ;
        RECT 286.520 0.820 286.800 1.100 ;
        RECT 287.440 0.820 287.720 1.100 ;
        RECT 288.100 0.820 288.380 1.100 ;
        RECT 288.760 0.820 289.040 1.100 ;
        RECT 289.680 0.820 289.960 1.100 ;
        RECT 290.340 0.820 290.620 1.100 ;
        RECT 291.000 0.820 291.280 1.100 ;
        RECT 291.920 0.820 292.200 1.100 ;
        RECT 292.580 0.820 292.860 1.100 ;
        RECT 293.240 0.820 293.520 1.100 ;
        RECT 294.160 0.820 294.440 1.100 ;
        RECT 294.820 0.820 295.100 1.100 ;
        RECT 295.480 0.820 295.760 1.100 ;
        RECT 296.400 0.820 296.680 1.100 ;
        RECT 297.060 0.820 297.340 1.100 ;
        RECT 297.720 0.820 298.000 1.100 ;
        RECT 298.640 0.820 298.920 1.100 ;
        RECT 299.300 0.820 299.580 1.100 ;
        RECT 299.960 0.820 300.240 1.100 ;
        RECT 301.000 0.820 301.280 1.100 ;
        RECT 302.000 0.820 302.280 1.100 ;
        RECT 302.660 0.820 302.940 1.100 ;
        RECT 303.320 0.820 303.600 1.100 ;
        RECT 304.240 0.820 304.520 1.100 ;
        RECT 304.900 0.820 305.180 1.100 ;
        RECT 305.560 0.820 305.840 1.100 ;
        RECT 306.480 0.820 306.760 1.100 ;
        RECT 307.140 0.820 307.420 1.100 ;
        RECT 307.800 0.820 308.080 1.100 ;
        RECT 308.720 0.820 309.000 1.100 ;
        RECT 309.380 0.820 309.660 1.100 ;
        RECT 310.040 0.820 310.320 1.100 ;
        RECT 310.800 0.820 311.080 1.100 ;
        RECT 312.120 0.820 312.400 1.100 ;
        RECT 314.320 0.820 314.600 1.100 ;
        RECT 314.980 0.820 315.260 1.100 ;
        RECT 315.640 0.820 315.920 1.100 ;
        RECT 316.560 0.820 316.840 1.100 ;
        RECT 317.220 0.820 317.500 1.100 ;
        RECT 317.880 0.820 318.160 1.100 ;
        RECT 318.800 0.820 319.080 1.100 ;
        RECT 319.460 0.820 319.740 1.100 ;
        RECT 320.120 0.820 320.400 1.100 ;
        RECT 321.160 0.820 321.440 1.100 ;
        RECT 322.160 0.820 322.440 1.100 ;
        RECT 322.820 0.820 323.100 1.100 ;
        RECT 323.480 0.820 323.760 1.100 ;
        RECT 324.400 0.820 324.680 1.100 ;
        RECT 325.060 0.820 325.340 1.100 ;
        RECT 325.720 0.820 326.000 1.100 ;
        RECT 326.640 0.820 326.920 1.100 ;
        RECT 327.300 0.820 327.580 1.100 ;
        RECT 327.960 0.820 328.240 1.100 ;
        RECT 328.880 0.820 329.160 1.100 ;
        RECT 329.540 0.820 329.820 1.100 ;
        RECT 330.200 0.820 330.480 1.100 ;
        RECT 331.120 0.820 331.400 1.100 ;
        RECT 331.780 0.820 332.060 1.100 ;
        RECT 332.440 0.820 332.720 1.100 ;
        RECT 333.360 0.820 333.640 1.100 ;
        RECT 334.020 0.820 334.300 1.100 ;
        RECT 334.680 0.820 334.960 1.100 ;
        RECT 335.600 0.820 335.880 1.100 ;
        RECT 336.260 0.820 336.540 1.100 ;
        RECT 336.920 0.820 337.200 1.100 ;
        RECT 337.840 0.820 338.120 1.100 ;
        RECT 338.500 0.820 338.780 1.100 ;
        RECT 339.160 0.820 339.440 1.100 ;
        RECT 340.080 0.820 340.360 1.100 ;
        RECT 340.740 0.820 341.020 1.100 ;
        RECT 341.400 0.820 341.680 1.100 ;
        RECT 342.440 0.820 342.720 1.100 ;
        RECT 343.440 0.820 343.720 1.100 ;
        RECT 344.100 0.820 344.380 1.100 ;
        RECT 344.760 0.820 345.040 1.100 ;
        RECT 345.680 0.820 345.960 1.100 ;
        RECT 346.340 0.820 346.620 1.100 ;
        RECT 347.000 0.820 347.280 1.100 ;
        RECT 347.920 0.820 348.200 1.100 ;
        RECT 348.580 0.820 348.860 1.100 ;
        RECT 349.240 0.820 349.520 1.100 ;
        RECT 350.160 0.820 350.440 1.100 ;
        RECT 350.820 0.820 351.100 1.100 ;
        RECT 351.480 0.820 351.760 1.100 ;
        RECT 352.240 0.820 352.520 1.100 ;
        RECT 353.560 0.820 353.840 1.100 ;
        RECT 355.760 0.820 356.040 1.100 ;
        RECT 356.420 0.820 356.700 1.100 ;
        RECT 357.080 0.820 357.360 1.100 ;
        RECT 358.000 0.820 358.280 1.100 ;
        RECT 358.660 0.820 358.940 1.100 ;
        RECT 359.320 0.820 359.600 1.100 ;
        RECT 360.240 0.820 360.520 1.100 ;
        RECT 360.900 0.820 361.180 1.100 ;
        RECT 361.560 0.820 361.840 1.100 ;
        RECT 362.600 0.820 362.880 1.100 ;
        RECT 363.600 0.820 363.880 1.100 ;
        RECT 364.260 0.820 364.540 1.100 ;
        RECT 364.920 0.820 365.200 1.100 ;
        RECT 365.840 0.820 366.120 1.100 ;
        RECT 366.500 0.820 366.780 1.100 ;
        RECT 367.160 0.820 367.440 1.100 ;
        RECT 368.080 0.820 368.360 1.100 ;
        RECT 368.740 0.820 369.020 1.100 ;
        RECT 369.400 0.820 369.680 1.100 ;
        RECT 370.320 0.820 370.600 1.100 ;
        RECT 370.980 0.820 371.260 1.100 ;
        RECT 371.640 0.820 371.920 1.100 ;
        RECT 372.560 0.820 372.840 1.100 ;
        RECT 373.220 0.820 373.500 1.100 ;
        RECT 373.880 0.820 374.160 1.100 ;
        RECT 374.800 0.820 375.080 1.100 ;
        RECT 375.460 0.820 375.740 1.100 ;
        RECT 376.120 0.820 376.400 1.100 ;
        RECT 377.040 0.820 377.320 1.100 ;
        RECT 377.700 0.820 377.980 1.100 ;
        RECT 378.360 0.820 378.640 1.100 ;
        RECT 379.280 0.820 379.560 1.100 ;
        RECT 379.940 0.820 380.220 1.100 ;
        RECT 380.600 0.820 380.880 1.100 ;
        RECT 381.520 0.820 381.800 1.100 ;
        RECT 382.180 0.820 382.460 1.100 ;
        RECT 382.840 0.820 383.120 1.100 ;
        RECT 383.880 0.820 384.160 1.100 ;
        RECT 384.880 0.820 385.160 1.100 ;
        RECT 385.540 0.820 385.820 1.100 ;
        RECT 386.200 0.820 386.480 1.100 ;
        RECT 387.120 0.820 387.400 1.100 ;
        RECT 387.780 0.820 388.060 1.100 ;
        RECT 388.440 0.820 388.720 1.100 ;
        RECT 389.360 0.820 389.640 1.100 ;
        RECT 390.020 0.820 390.300 1.100 ;
        RECT 390.680 0.820 390.960 1.100 ;
        RECT 391.600 0.820 391.880 1.100 ;
        RECT 392.260 0.820 392.540 1.100 ;
        RECT 392.920 0.820 393.200 1.100 ;
        RECT 393.840 0.820 394.120 1.100 ;
        RECT 394.500 0.820 394.780 1.100 ;
        RECT 395.160 0.820 395.440 1.100 ;
        RECT 395.920 0.820 396.200 1.100 ;
        RECT 397.240 0.820 397.520 1.100 ;
        RECT 399.440 0.820 399.720 1.100 ;
        RECT 400.100 0.820 400.380 1.100 ;
        RECT 400.760 0.820 401.040 1.100 ;
        RECT 401.680 0.820 401.960 1.100 ;
        RECT 402.340 0.820 402.620 1.100 ;
        RECT 403.000 0.820 403.280 1.100 ;
        RECT 404.040 0.820 404.320 1.100 ;
        RECT 405.040 0.820 405.320 1.100 ;
        RECT 405.700 0.820 405.980 1.100 ;
        RECT 406.360 0.820 406.640 1.100 ;
        RECT 407.280 0.820 407.560 1.100 ;
        RECT 407.940 0.820 408.220 1.100 ;
        RECT 408.600 0.820 408.880 1.100 ;
        RECT 409.520 0.820 409.800 1.100 ;
        RECT 410.180 0.820 410.460 1.100 ;
        RECT 410.840 0.820 411.120 1.100 ;
        RECT 411.760 0.820 412.040 1.100 ;
        RECT 412.420 0.820 412.700 1.100 ;
        RECT 413.080 0.820 413.360 1.100 ;
        RECT 414.000 0.820 414.280 1.100 ;
        RECT 414.660 0.820 414.940 1.100 ;
        RECT 415.320 0.820 415.600 1.100 ;
        RECT 416.240 0.820 416.520 1.100 ;
        RECT 416.900 0.820 417.180 1.100 ;
        RECT 417.560 0.820 417.840 1.100 ;
        RECT 418.480 0.820 418.760 1.100 ;
        RECT 419.140 0.820 419.420 1.100 ;
        RECT 419.800 0.820 420.080 1.100 ;
        RECT 420.720 0.820 421.000 1.100 ;
        RECT 421.380 0.820 421.660 1.100 ;
        RECT 422.040 0.820 422.320 1.100 ;
        RECT 422.960 0.820 423.240 1.100 ;
        RECT 423.620 0.820 423.900 1.100 ;
        RECT 424.280 0.820 424.560 1.100 ;
        RECT 425.320 0.820 425.600 1.100 ;
        RECT 426.320 0.820 426.600 1.100 ;
        RECT 426.980 0.820 427.260 1.100 ;
        RECT 427.640 0.820 427.920 1.100 ;
        RECT 428.560 0.820 428.840 1.100 ;
        RECT 429.220 0.820 429.500 1.100 ;
        RECT 429.880 0.820 430.160 1.100 ;
        RECT 430.800 0.820 431.080 1.100 ;
        RECT 431.460 0.820 431.740 1.100 ;
        RECT 432.120 0.820 432.400 1.100 ;
        RECT 433.040 0.820 433.320 1.100 ;
        RECT 433.700 0.820 433.980 1.100 ;
        RECT 434.360 0.820 434.640 1.100 ;
        RECT 435.280 0.820 435.560 1.100 ;
        RECT 435.940 0.820 436.220 1.100 ;
        RECT 436.600 0.820 436.880 1.100 ;
        RECT 437.360 0.820 437.640 1.100 ;
        RECT 438.680 0.820 438.960 1.100 ;
        RECT 440.880 0.820 441.160 1.100 ;
        RECT 441.540 0.820 441.820 1.100 ;
        RECT 442.200 0.820 442.480 1.100 ;
        RECT 443.120 0.820 443.400 1.100 ;
        RECT 443.780 0.820 444.060 1.100 ;
        RECT 444.440 0.820 444.720 1.100 ;
        RECT 445.480 0.820 445.760 1.100 ;
        RECT 446.480 0.820 446.760 1.100 ;
        RECT 447.140 0.820 447.420 1.100 ;
        RECT 447.800 0.820 448.080 1.100 ;
        RECT 448.720 0.820 449.000 1.100 ;
        RECT 449.380 0.820 449.660 1.100 ;
        RECT 450.040 0.820 450.320 1.100 ;
        RECT 450.960 0.820 451.240 1.100 ;
        RECT 451.620 0.820 451.900 1.100 ;
        RECT 452.280 0.820 452.560 1.100 ;
        RECT 453.200 0.820 453.480 1.100 ;
        RECT 453.860 0.820 454.140 1.100 ;
        RECT 454.520 0.820 454.800 1.100 ;
        RECT 455.440 0.820 455.720 1.100 ;
        RECT 456.100 0.820 456.380 1.100 ;
        RECT 456.760 0.820 457.040 1.100 ;
        RECT 457.680 0.820 457.960 1.100 ;
        RECT 458.340 0.820 458.620 1.100 ;
        RECT 459.000 0.820 459.280 1.100 ;
        RECT 459.920 0.820 460.200 1.100 ;
        RECT 460.580 0.820 460.860 1.100 ;
        RECT 461.240 0.820 461.520 1.100 ;
        RECT 462.160 0.820 462.440 1.100 ;
        RECT 462.820 0.820 463.100 1.100 ;
        RECT 463.480 0.820 463.760 1.100 ;
        RECT 464.400 0.820 464.680 1.100 ;
        RECT 465.060 0.820 465.340 1.100 ;
        RECT 465.720 0.820 466.000 1.100 ;
        RECT 466.760 0.820 467.040 1.100 ;
        RECT 467.760 0.820 468.040 1.100 ;
        RECT 468.420 0.820 468.700 1.100 ;
        RECT 469.080 0.820 469.360 1.100 ;
        RECT 470.000 0.820 470.280 1.100 ;
        RECT 470.660 0.820 470.940 1.100 ;
        RECT 471.320 0.820 471.600 1.100 ;
        RECT 472.240 0.820 472.520 1.100 ;
        RECT 472.900 0.820 473.180 1.100 ;
        RECT 473.560 0.820 473.840 1.100 ;
        RECT 474.480 0.820 474.760 1.100 ;
        RECT 475.140 0.820 475.420 1.100 ;
        RECT 475.800 0.820 476.080 1.100 ;
        RECT 476.720 0.820 477.000 1.100 ;
        RECT 477.380 0.820 477.660 1.100 ;
        RECT 478.040 0.820 478.320 1.100 ;
        RECT 478.960 0.820 479.240 1.100 ;
        RECT 479.620 0.820 479.900 1.100 ;
        RECT 480.280 0.820 480.560 1.100 ;
        RECT 481.040 0.820 481.320 1.100 ;
        RECT 482.360 0.820 482.640 1.100 ;
        RECT 484.560 0.820 484.840 1.100 ;
        RECT 485.220 0.820 485.500 1.100 ;
        RECT 485.880 0.820 486.160 1.100 ;
        RECT 486.920 0.820 487.200 1.100 ;
        RECT 487.920 0.820 488.200 1.100 ;
        RECT 488.580 0.820 488.860 1.100 ;
        RECT 489.240 0.820 489.520 1.100 ;
        RECT 490.160 0.820 490.440 1.100 ;
        RECT 490.820 0.820 491.100 1.100 ;
        RECT 491.480 0.820 491.760 1.100 ;
        RECT 492.400 0.820 492.680 1.100 ;
        RECT 493.060 0.820 493.340 1.100 ;
        RECT 493.720 0.820 494.000 1.100 ;
        RECT 494.640 0.820 494.920 1.100 ;
        RECT 495.300 0.820 495.580 1.100 ;
        RECT 495.960 0.820 496.240 1.100 ;
        RECT 496.880 0.820 497.160 1.100 ;
        RECT 497.540 0.820 497.820 1.100 ;
        RECT 498.200 0.820 498.480 1.100 ;
        RECT 499.120 0.820 499.400 1.100 ;
        RECT 499.780 0.820 500.060 1.100 ;
        RECT 500.440 0.820 500.720 1.100 ;
        RECT 501.360 0.820 501.640 1.100 ;
        RECT 502.020 0.820 502.300 1.100 ;
        RECT 502.680 0.820 502.960 1.100 ;
        RECT 503.600 0.820 503.880 1.100 ;
        RECT 504.260 0.820 504.540 1.100 ;
        RECT 504.920 0.820 505.200 1.100 ;
        RECT 505.840 0.820 506.120 1.100 ;
        RECT 506.500 0.820 506.780 1.100 ;
        RECT 507.160 0.820 507.440 1.100 ;
        RECT 508.200 0.820 508.480 1.100 ;
        RECT 509.200 0.820 509.480 1.100 ;
        RECT 509.860 0.820 510.140 1.100 ;
        RECT 510.520 0.820 510.800 1.100 ;
        RECT 511.440 0.820 511.720 1.100 ;
        RECT 512.100 0.820 512.380 1.100 ;
        RECT 512.760 0.820 513.040 1.100 ;
        RECT 513.680 0.820 513.960 1.100 ;
        RECT 514.340 0.820 514.620 1.100 ;
        RECT 515.000 0.820 515.280 1.100 ;
        RECT 515.920 0.820 516.200 1.100 ;
        RECT 516.580 0.820 516.860 1.100 ;
        RECT 517.240 0.820 517.520 1.100 ;
        RECT 518.160 0.820 518.440 1.100 ;
        RECT 518.820 0.820 519.100 1.100 ;
        RECT 519.480 0.820 519.760 1.100 ;
        RECT 520.400 0.820 520.680 1.100 ;
        RECT 521.060 0.820 521.340 1.100 ;
        RECT 521.720 0.820 522.000 1.100 ;
        RECT 522.480 0.820 522.760 1.100 ;
        RECT 523.800 0.820 524.080 1.100 ;
        RECT 526.000 0.820 526.280 1.100 ;
        RECT 526.660 0.820 526.940 1.100 ;
        RECT 527.320 0.820 527.600 1.100 ;
        RECT 528.360 0.820 528.640 1.100 ;
        RECT 529.360 0.820 529.640 1.100 ;
        RECT 530.020 0.820 530.300 1.100 ;
        RECT 530.680 0.820 530.960 1.100 ;
        RECT 531.600 0.820 531.880 1.100 ;
        RECT 532.260 0.820 532.540 1.100 ;
        RECT 532.920 0.820 533.200 1.100 ;
        RECT 533.840 0.820 534.120 1.100 ;
        RECT 534.500 0.820 534.780 1.100 ;
        RECT 535.160 0.820 535.440 1.100 ;
        RECT 536.080 0.820 536.360 1.100 ;
        RECT 536.740 0.820 537.020 1.100 ;
        RECT 537.400 0.820 537.680 1.100 ;
        RECT 538.320 0.820 538.600 1.100 ;
        RECT 538.980 0.820 539.260 1.100 ;
        RECT 539.640 0.820 539.920 1.100 ;
        RECT 540.560 0.820 540.840 1.100 ;
        RECT 541.220 0.820 541.500 1.100 ;
        RECT 541.880 0.820 542.160 1.100 ;
        RECT 542.800 0.820 543.080 1.100 ;
        RECT 543.460 0.820 543.740 1.100 ;
        RECT 544.120 0.820 544.400 1.100 ;
        RECT 545.040 0.820 545.320 1.100 ;
        RECT 545.700 0.820 545.980 1.100 ;
        RECT 546.360 0.820 546.640 1.100 ;
        RECT 547.280 0.820 547.560 1.100 ;
        RECT 547.940 0.820 548.220 1.100 ;
        RECT 548.600 0.820 548.880 1.100 ;
        RECT 549.640 0.820 549.920 1.100 ;
        RECT 550.640 0.820 550.920 1.100 ;
        RECT 551.300 0.820 551.580 1.100 ;
        RECT 551.960 0.820 552.240 1.100 ;
        RECT 552.880 0.820 553.160 1.100 ;
        RECT 553.540 0.820 553.820 1.100 ;
        RECT 554.200 0.820 554.480 1.100 ;
        RECT 555.120 0.820 555.400 1.100 ;
        RECT 555.780 0.820 556.060 1.100 ;
        RECT 556.440 0.820 556.720 1.100 ;
        RECT 557.360 0.820 557.640 1.100 ;
        RECT 558.020 0.820 558.300 1.100 ;
        RECT 558.680 0.820 558.960 1.100 ;
        RECT 559.600 0.820 559.880 1.100 ;
        RECT 560.260 0.820 560.540 1.100 ;
        RECT 560.920 0.820 561.200 1.100 ;
        RECT 561.840 0.820 562.120 1.100 ;
        RECT 562.500 0.820 562.780 1.100 ;
        RECT 563.160 0.820 563.440 1.100 ;
        RECT 564.080 0.820 564.360 1.100 ;
        RECT 564.740 0.820 565.020 1.100 ;
        RECT 565.400 0.820 565.680 1.100 ;
        RECT 566.160 0.820 566.440 1.100 ;
        RECT 567.480 0.820 567.760 1.100 ;
        RECT 569.800 0.820 570.080 1.100 ;
        RECT 570.800 0.820 571.080 1.100 ;
        RECT 571.460 0.820 571.740 1.100 ;
        RECT 572.120 0.820 572.400 1.100 ;
        RECT 573.040 0.820 573.320 1.100 ;
        RECT 573.700 0.820 573.980 1.100 ;
        RECT 574.360 0.820 574.640 1.100 ;
        RECT 575.280 0.820 575.560 1.100 ;
        RECT 575.940 0.820 576.220 1.100 ;
        RECT 576.600 0.820 576.880 1.100 ;
        RECT 577.520 0.820 577.800 1.100 ;
        RECT 578.180 0.820 578.460 1.100 ;
        RECT 578.840 0.820 579.120 1.100 ;
        RECT 579.760 0.820 580.040 1.100 ;
        RECT 580.420 0.820 580.700 1.100 ;
        RECT 581.080 0.820 581.360 1.100 ;
        RECT 582.000 0.820 582.280 1.100 ;
        RECT 582.660 0.820 582.940 1.100 ;
        RECT 583.320 0.820 583.600 1.100 ;
        RECT 584.240 0.820 584.520 1.100 ;
        RECT 584.900 0.820 585.180 1.100 ;
        RECT 585.560 0.820 585.840 1.100 ;
        RECT 586.480 0.820 586.760 1.100 ;
        RECT 587.140 0.820 587.420 1.100 ;
        RECT 587.800 0.820 588.080 1.100 ;
        RECT 588.720 0.820 589.000 1.100 ;
        RECT 589.380 0.820 589.660 1.100 ;
        RECT 590.040 0.820 590.320 1.100 ;
        RECT 591.080 0.820 591.360 1.100 ;
        RECT 592.080 0.820 592.360 1.100 ;
        RECT 592.740 0.820 593.020 1.100 ;
        RECT 593.400 0.820 593.680 1.100 ;
        RECT 594.320 0.820 594.600 1.100 ;
        RECT 594.980 0.820 595.260 1.100 ;
        RECT 595.640 0.820 595.920 1.100 ;
        RECT 596.560 0.820 596.840 1.100 ;
        RECT 597.220 0.820 597.500 1.100 ;
        RECT 597.880 0.820 598.160 1.100 ;
        RECT 598.800 0.820 599.080 1.100 ;
        RECT 599.460 0.820 599.740 1.100 ;
        RECT 600.120 0.820 600.400 1.100 ;
        RECT 601.040 0.820 601.320 1.100 ;
        RECT 601.700 0.820 601.980 1.100 ;
        RECT 602.360 0.820 602.640 1.100 ;
        RECT 603.280 0.820 603.560 1.100 ;
        RECT 603.940 0.820 604.220 1.100 ;
        RECT 604.600 0.820 604.880 1.100 ;
        RECT 605.520 0.820 605.800 1.100 ;
        RECT 606.180 0.820 606.460 1.100 ;
        RECT 606.840 0.820 607.120 1.100 ;
        RECT 607.600 0.820 607.880 1.100 ;
        RECT 608.920 0.820 609.200 1.100 ;
        RECT 611.240 0.820 611.520 1.100 ;
        RECT 612.240 0.820 612.520 1.100 ;
        RECT 612.900 0.820 613.180 1.100 ;
        RECT 613.560 0.820 613.840 1.100 ;
        RECT 614.480 0.820 614.760 1.100 ;
        RECT 615.140 0.820 615.420 1.100 ;
        RECT 615.800 0.820 616.080 1.100 ;
        RECT 616.720 0.820 617.000 1.100 ;
        RECT 617.380 0.820 617.660 1.100 ;
        RECT 618.040 0.820 618.320 1.100 ;
        RECT 618.960 0.820 619.240 1.100 ;
        RECT 619.620 0.820 619.900 1.100 ;
        RECT 620.280 0.820 620.560 1.100 ;
        RECT 621.200 0.820 621.480 1.100 ;
        RECT 621.860 0.820 622.140 1.100 ;
        RECT 622.520 0.820 622.800 1.100 ;
        RECT 623.440 0.820 623.720 1.100 ;
        RECT 624.100 0.820 624.380 1.100 ;
        RECT 624.760 0.820 625.040 1.100 ;
        RECT 625.680 0.820 625.960 1.100 ;
        RECT 626.340 0.820 626.620 1.100 ;
        RECT 627.000 0.820 627.280 1.100 ;
        RECT 627.920 0.820 628.200 1.100 ;
        RECT 628.580 0.820 628.860 1.100 ;
        RECT 629.240 0.820 629.520 1.100 ;
        RECT 630.160 0.820 630.440 1.100 ;
        RECT 630.820 0.820 631.100 1.100 ;
        RECT 631.480 0.820 631.760 1.100 ;
        RECT 632.520 0.820 632.800 1.100 ;
        RECT 633.520 0.820 633.800 1.100 ;
        RECT 634.180 0.820 634.460 1.100 ;
        RECT 634.840 0.820 635.120 1.100 ;
        RECT 635.760 0.820 636.040 1.100 ;
        RECT 636.420 0.820 636.700 1.100 ;
        RECT 637.080 0.820 637.360 1.100 ;
        RECT 638.000 0.820 638.280 1.100 ;
        RECT 638.660 0.820 638.940 1.100 ;
        RECT 639.320 0.820 639.600 1.100 ;
        RECT 640.240 0.820 640.520 1.100 ;
        RECT 640.900 0.820 641.180 1.100 ;
        RECT 641.560 0.820 641.840 1.100 ;
        RECT 642.480 0.820 642.760 1.100 ;
        RECT 643.140 0.820 643.420 1.100 ;
        RECT 643.800 0.820 644.080 1.100 ;
        RECT 644.720 0.820 645.000 1.100 ;
        RECT 645.380 0.820 645.660 1.100 ;
        RECT 646.040 0.820 646.320 1.100 ;
        RECT 646.960 0.820 647.240 1.100 ;
        RECT 647.620 0.820 647.900 1.100 ;
        RECT 648.280 0.820 648.560 1.100 ;
        RECT 649.200 0.820 649.480 1.100 ;
        RECT 649.860 0.820 650.140 1.100 ;
        RECT 650.520 0.820 650.800 1.100 ;
        RECT 651.280 0.820 651.560 1.100 ;
        RECT 652.600 0.820 652.880 1.100 ;
        RECT 654.920 0.820 655.200 1.100 ;
        RECT 655.920 0.820 656.200 1.100 ;
        RECT 656.580 0.820 656.860 1.100 ;
        RECT 657.240 0.820 657.520 1.100 ;
        RECT 658.160 0.820 658.440 1.100 ;
        RECT 658.820 0.820 659.100 1.100 ;
        RECT 659.480 0.820 659.760 1.100 ;
        RECT 660.400 0.820 660.680 1.100 ;
        RECT 661.060 0.820 661.340 1.100 ;
        RECT 661.720 0.820 662.000 1.100 ;
        RECT 662.640 0.820 662.920 1.100 ;
        RECT 663.300 0.820 663.580 1.100 ;
        RECT 663.960 0.820 664.240 1.100 ;
        RECT 664.880 0.820 665.160 1.100 ;
        RECT 665.540 0.820 665.820 1.100 ;
        RECT 666.200 0.820 666.480 1.100 ;
        RECT 667.120 0.820 667.400 1.100 ;
        RECT 667.780 0.820 668.060 1.100 ;
        RECT 668.440 0.820 668.720 1.100 ;
        RECT 669.360 0.820 669.640 1.100 ;
        RECT 670.020 0.820 670.300 1.100 ;
        RECT 670.680 0.820 670.960 1.100 ;
        RECT 671.600 0.820 671.880 1.100 ;
        RECT 672.260 0.820 672.540 1.100 ;
        RECT 672.920 0.820 673.200 1.100 ;
        RECT 673.840 0.820 674.120 1.100 ;
        RECT 674.500 0.820 674.780 1.100 ;
        RECT 675.160 0.820 675.440 1.100 ;
        RECT 676.200 0.820 676.480 1.100 ;
        RECT 677.200 0.820 677.480 1.100 ;
        RECT 677.860 0.820 678.140 1.100 ;
        RECT 678.520 0.820 678.800 1.100 ;
        RECT 679.540 0.820 679.820 1.100 ;
      LAYER Metal3 ;
        RECT 0.765 58.745 1.145 59.125 ;
        RECT 11.055 58.745 11.435 59.125 ;
        RECT 21.340 58.745 21.720 59.125 ;
        RECT 31.630 58.745 32.010 59.125 ;
        RECT 41.915 58.745 42.295 59.125 ;
        RECT 43.335 58.745 43.715 59.125 ;
        RECT 53.625 58.745 54.005 59.125 ;
        RECT 63.910 58.745 64.290 59.125 ;
        RECT 74.200 58.745 74.580 59.125 ;
        RECT 84.485 58.745 84.865 59.125 ;
        RECT 85.905 58.745 86.285 59.125 ;
        RECT 96.195 58.745 96.575 59.125 ;
        RECT 106.480 58.745 106.860 59.125 ;
        RECT 116.770 58.745 117.150 59.125 ;
        RECT 127.055 58.745 127.435 59.125 ;
        RECT 128.475 58.745 128.855 59.125 ;
        RECT 138.765 58.745 139.145 59.125 ;
        RECT 149.050 58.745 149.430 59.125 ;
        RECT 159.340 58.745 159.720 59.125 ;
        RECT 169.625 58.745 170.005 59.125 ;
        RECT 171.045 58.745 171.425 59.125 ;
        RECT 181.335 58.745 181.715 59.125 ;
        RECT 191.620 58.745 192.000 59.125 ;
        RECT 201.910 58.745 202.290 59.125 ;
        RECT 212.195 58.745 212.575 59.125 ;
        RECT 213.615 58.745 213.995 59.125 ;
        RECT 223.905 58.745 224.285 59.125 ;
        RECT 234.190 58.745 234.570 59.125 ;
        RECT 244.480 58.745 244.860 59.125 ;
        RECT 254.765 58.745 255.145 59.125 ;
        RECT 256.185 58.745 256.565 59.125 ;
        RECT 266.475 58.745 266.855 59.125 ;
        RECT 276.760 58.745 277.140 59.125 ;
        RECT 287.050 58.745 287.430 59.125 ;
        RECT 297.335 58.745 297.715 59.125 ;
        RECT 298.755 58.745 299.135 59.125 ;
        RECT 309.045 58.745 309.425 59.125 ;
        RECT 319.330 58.745 319.710 59.125 ;
        RECT 329.620 58.745 330.000 59.125 ;
        RECT 339.905 58.745 340.285 59.125 ;
        RECT 341.325 58.745 341.705 59.125 ;
        RECT 351.615 58.745 351.995 59.125 ;
        RECT 361.900 58.745 362.280 59.125 ;
        RECT 372.190 58.745 372.570 59.125 ;
        RECT 382.475 58.745 382.855 59.125 ;
        RECT 383.895 58.745 384.275 59.125 ;
        RECT 394.185 58.745 394.565 59.125 ;
        RECT 404.470 58.745 404.850 59.125 ;
        RECT 414.760 58.745 415.140 59.125 ;
        RECT 425.045 58.745 425.425 59.125 ;
        RECT 426.465 58.745 426.845 59.125 ;
        RECT 436.755 58.745 437.135 59.125 ;
        RECT 447.040 58.745 447.420 59.125 ;
        RECT 457.330 58.745 457.710 59.125 ;
        RECT 467.615 58.745 467.995 59.125 ;
        RECT 469.035 58.745 469.415 59.125 ;
        RECT 479.325 58.745 479.705 59.125 ;
        RECT 489.610 58.745 489.990 59.125 ;
        RECT 499.900 58.745 500.280 59.125 ;
        RECT 510.185 58.745 510.565 59.125 ;
        RECT 511.605 58.745 511.985 59.125 ;
        RECT 521.895 58.745 522.275 59.125 ;
        RECT 532.180 58.745 532.560 59.125 ;
        RECT 542.470 58.745 542.850 59.125 ;
        RECT 552.755 58.745 553.135 59.125 ;
        RECT 554.175 58.745 554.555 59.125 ;
        RECT 564.465 58.745 564.845 59.125 ;
        RECT 574.750 58.745 575.130 59.125 ;
        RECT 585.040 58.745 585.420 59.125 ;
        RECT 595.325 58.745 595.705 59.125 ;
        RECT 596.745 58.745 597.125 59.125 ;
        RECT 607.035 58.745 607.415 59.125 ;
        RECT 617.320 58.745 617.700 59.125 ;
        RECT 627.610 58.745 627.990 59.125 ;
        RECT 637.895 58.745 638.275 59.125 ;
        RECT 639.315 58.745 639.695 59.125 ;
        RECT 649.605 58.745 649.985 59.125 ;
        RECT 659.890 58.745 660.270 59.125 ;
        RECT 670.180 58.745 670.560 59.125 ;
        RECT 680.465 58.745 680.845 59.125 ;
        RECT 0.765 58.085 1.145 58.465 ;
        RECT 11.055 58.085 11.435 58.465 ;
        RECT 21.340 58.085 21.720 58.465 ;
        RECT 31.630 58.085 32.010 58.465 ;
        RECT 41.915 58.085 42.295 58.465 ;
        RECT 43.335 58.085 43.715 58.465 ;
        RECT 53.625 58.085 54.005 58.465 ;
        RECT 63.910 58.085 64.290 58.465 ;
        RECT 74.200 58.085 74.580 58.465 ;
        RECT 84.485 58.085 84.865 58.465 ;
        RECT 85.905 58.085 86.285 58.465 ;
        RECT 96.195 58.085 96.575 58.465 ;
        RECT 106.480 58.085 106.860 58.465 ;
        RECT 116.770 58.085 117.150 58.465 ;
        RECT 127.055 58.085 127.435 58.465 ;
        RECT 128.475 58.085 128.855 58.465 ;
        RECT 138.765 58.085 139.145 58.465 ;
        RECT 149.050 58.085 149.430 58.465 ;
        RECT 159.340 58.085 159.720 58.465 ;
        RECT 169.625 58.085 170.005 58.465 ;
        RECT 171.045 58.085 171.425 58.465 ;
        RECT 181.335 58.085 181.715 58.465 ;
        RECT 191.620 58.085 192.000 58.465 ;
        RECT 201.910 58.085 202.290 58.465 ;
        RECT 212.195 58.085 212.575 58.465 ;
        RECT 213.615 58.085 213.995 58.465 ;
        RECT 223.905 58.085 224.285 58.465 ;
        RECT 234.190 58.085 234.570 58.465 ;
        RECT 244.480 58.085 244.860 58.465 ;
        RECT 254.765 58.085 255.145 58.465 ;
        RECT 256.185 58.085 256.565 58.465 ;
        RECT 266.475 58.085 266.855 58.465 ;
        RECT 276.760 58.085 277.140 58.465 ;
        RECT 287.050 58.085 287.430 58.465 ;
        RECT 297.335 58.085 297.715 58.465 ;
        RECT 298.755 58.085 299.135 58.465 ;
        RECT 309.045 58.085 309.425 58.465 ;
        RECT 319.330 58.085 319.710 58.465 ;
        RECT 329.620 58.085 330.000 58.465 ;
        RECT 339.905 58.085 340.285 58.465 ;
        RECT 341.325 58.085 341.705 58.465 ;
        RECT 351.615 58.085 351.995 58.465 ;
        RECT 361.900 58.085 362.280 58.465 ;
        RECT 372.190 58.085 372.570 58.465 ;
        RECT 382.475 58.085 382.855 58.465 ;
        RECT 383.895 58.085 384.275 58.465 ;
        RECT 394.185 58.085 394.565 58.465 ;
        RECT 404.470 58.085 404.850 58.465 ;
        RECT 414.760 58.085 415.140 58.465 ;
        RECT 425.045 58.085 425.425 58.465 ;
        RECT 426.465 58.085 426.845 58.465 ;
        RECT 436.755 58.085 437.135 58.465 ;
        RECT 447.040 58.085 447.420 58.465 ;
        RECT 457.330 58.085 457.710 58.465 ;
        RECT 467.615 58.085 467.995 58.465 ;
        RECT 469.035 58.085 469.415 58.465 ;
        RECT 479.325 58.085 479.705 58.465 ;
        RECT 489.610 58.085 489.990 58.465 ;
        RECT 499.900 58.085 500.280 58.465 ;
        RECT 510.185 58.085 510.565 58.465 ;
        RECT 511.605 58.085 511.985 58.465 ;
        RECT 521.895 58.085 522.275 58.465 ;
        RECT 532.180 58.085 532.560 58.465 ;
        RECT 542.470 58.085 542.850 58.465 ;
        RECT 552.755 58.085 553.135 58.465 ;
        RECT 554.175 58.085 554.555 58.465 ;
        RECT 564.465 58.085 564.845 58.465 ;
        RECT 574.750 58.085 575.130 58.465 ;
        RECT 585.040 58.085 585.420 58.465 ;
        RECT 595.325 58.085 595.705 58.465 ;
        RECT 596.745 58.085 597.125 58.465 ;
        RECT 607.035 58.085 607.415 58.465 ;
        RECT 617.320 58.085 617.700 58.465 ;
        RECT 627.610 58.085 627.990 58.465 ;
        RECT 637.895 58.085 638.275 58.465 ;
        RECT 639.315 58.085 639.695 58.465 ;
        RECT 649.605 58.085 649.985 58.465 ;
        RECT 659.890 58.085 660.270 58.465 ;
        RECT 670.180 58.085 670.560 58.465 ;
        RECT 680.465 58.085 680.845 58.465 ;
        RECT 0.765 57.425 1.145 57.805 ;
        RECT 11.055 57.425 11.435 57.805 ;
        RECT 21.340 57.425 21.720 57.805 ;
        RECT 31.630 57.425 32.010 57.805 ;
        RECT 41.915 57.425 42.295 57.805 ;
        RECT 43.335 57.425 43.715 57.805 ;
        RECT 53.625 57.425 54.005 57.805 ;
        RECT 63.910 57.425 64.290 57.805 ;
        RECT 74.200 57.425 74.580 57.805 ;
        RECT 84.485 57.425 84.865 57.805 ;
        RECT 85.905 57.425 86.285 57.805 ;
        RECT 96.195 57.425 96.575 57.805 ;
        RECT 106.480 57.425 106.860 57.805 ;
        RECT 116.770 57.425 117.150 57.805 ;
        RECT 127.055 57.425 127.435 57.805 ;
        RECT 128.475 57.425 128.855 57.805 ;
        RECT 138.765 57.425 139.145 57.805 ;
        RECT 149.050 57.425 149.430 57.805 ;
        RECT 159.340 57.425 159.720 57.805 ;
        RECT 169.625 57.425 170.005 57.805 ;
        RECT 171.045 57.425 171.425 57.805 ;
        RECT 181.335 57.425 181.715 57.805 ;
        RECT 191.620 57.425 192.000 57.805 ;
        RECT 201.910 57.425 202.290 57.805 ;
        RECT 212.195 57.425 212.575 57.805 ;
        RECT 213.615 57.425 213.995 57.805 ;
        RECT 223.905 57.425 224.285 57.805 ;
        RECT 234.190 57.425 234.570 57.805 ;
        RECT 244.480 57.425 244.860 57.805 ;
        RECT 254.765 57.425 255.145 57.805 ;
        RECT 256.185 57.425 256.565 57.805 ;
        RECT 266.475 57.425 266.855 57.805 ;
        RECT 276.760 57.425 277.140 57.805 ;
        RECT 287.050 57.425 287.430 57.805 ;
        RECT 297.335 57.425 297.715 57.805 ;
        RECT 298.755 57.425 299.135 57.805 ;
        RECT 309.045 57.425 309.425 57.805 ;
        RECT 319.330 57.425 319.710 57.805 ;
        RECT 329.620 57.425 330.000 57.805 ;
        RECT 339.905 57.425 340.285 57.805 ;
        RECT 341.325 57.425 341.705 57.805 ;
        RECT 351.615 57.425 351.995 57.805 ;
        RECT 361.900 57.425 362.280 57.805 ;
        RECT 372.190 57.425 372.570 57.805 ;
        RECT 382.475 57.425 382.855 57.805 ;
        RECT 383.895 57.425 384.275 57.805 ;
        RECT 394.185 57.425 394.565 57.805 ;
        RECT 404.470 57.425 404.850 57.805 ;
        RECT 414.760 57.425 415.140 57.805 ;
        RECT 425.045 57.425 425.425 57.805 ;
        RECT 426.465 57.425 426.845 57.805 ;
        RECT 436.755 57.425 437.135 57.805 ;
        RECT 447.040 57.425 447.420 57.805 ;
        RECT 457.330 57.425 457.710 57.805 ;
        RECT 467.615 57.425 467.995 57.805 ;
        RECT 469.035 57.425 469.415 57.805 ;
        RECT 479.325 57.425 479.705 57.805 ;
        RECT 489.610 57.425 489.990 57.805 ;
        RECT 499.900 57.425 500.280 57.805 ;
        RECT 510.185 57.425 510.565 57.805 ;
        RECT 511.605 57.425 511.985 57.805 ;
        RECT 521.895 57.425 522.275 57.805 ;
        RECT 532.180 57.425 532.560 57.805 ;
        RECT 542.470 57.425 542.850 57.805 ;
        RECT 552.755 57.425 553.135 57.805 ;
        RECT 554.175 57.425 554.555 57.805 ;
        RECT 564.465 57.425 564.845 57.805 ;
        RECT 574.750 57.425 575.130 57.805 ;
        RECT 585.040 57.425 585.420 57.805 ;
        RECT 595.325 57.425 595.705 57.805 ;
        RECT 596.745 57.425 597.125 57.805 ;
        RECT 607.035 57.425 607.415 57.805 ;
        RECT 617.320 57.425 617.700 57.805 ;
        RECT 627.610 57.425 627.990 57.805 ;
        RECT 637.895 57.425 638.275 57.805 ;
        RECT 639.315 57.425 639.695 57.805 ;
        RECT 649.605 57.425 649.985 57.805 ;
        RECT 659.890 57.425 660.270 57.805 ;
        RECT 670.180 57.425 670.560 57.805 ;
        RECT 680.465 57.425 680.845 57.805 ;
        RECT 0.765 56.765 1.145 57.145 ;
        RECT 11.055 56.765 11.435 57.145 ;
        RECT 21.340 56.765 21.720 57.145 ;
        RECT 31.630 56.765 32.010 57.145 ;
        RECT 41.915 56.765 42.295 57.145 ;
        RECT 43.335 56.765 43.715 57.145 ;
        RECT 53.625 56.765 54.005 57.145 ;
        RECT 63.910 56.765 64.290 57.145 ;
        RECT 74.200 56.765 74.580 57.145 ;
        RECT 84.485 56.765 84.865 57.145 ;
        RECT 85.905 56.765 86.285 57.145 ;
        RECT 96.195 56.765 96.575 57.145 ;
        RECT 106.480 56.765 106.860 57.145 ;
        RECT 116.770 56.765 117.150 57.145 ;
        RECT 127.055 56.765 127.435 57.145 ;
        RECT 128.475 56.765 128.855 57.145 ;
        RECT 138.765 56.765 139.145 57.145 ;
        RECT 149.050 56.765 149.430 57.145 ;
        RECT 159.340 56.765 159.720 57.145 ;
        RECT 169.625 56.765 170.005 57.145 ;
        RECT 171.045 56.765 171.425 57.145 ;
        RECT 181.335 56.765 181.715 57.145 ;
        RECT 191.620 56.765 192.000 57.145 ;
        RECT 201.910 56.765 202.290 57.145 ;
        RECT 212.195 56.765 212.575 57.145 ;
        RECT 213.615 56.765 213.995 57.145 ;
        RECT 223.905 56.765 224.285 57.145 ;
        RECT 234.190 56.765 234.570 57.145 ;
        RECT 244.480 56.765 244.860 57.145 ;
        RECT 254.765 56.765 255.145 57.145 ;
        RECT 256.185 56.765 256.565 57.145 ;
        RECT 266.475 56.765 266.855 57.145 ;
        RECT 276.760 56.765 277.140 57.145 ;
        RECT 287.050 56.765 287.430 57.145 ;
        RECT 297.335 56.765 297.715 57.145 ;
        RECT 298.755 56.765 299.135 57.145 ;
        RECT 309.045 56.765 309.425 57.145 ;
        RECT 319.330 56.765 319.710 57.145 ;
        RECT 329.620 56.765 330.000 57.145 ;
        RECT 339.905 56.765 340.285 57.145 ;
        RECT 341.325 56.765 341.705 57.145 ;
        RECT 351.615 56.765 351.995 57.145 ;
        RECT 361.900 56.765 362.280 57.145 ;
        RECT 372.190 56.765 372.570 57.145 ;
        RECT 382.475 56.765 382.855 57.145 ;
        RECT 383.895 56.765 384.275 57.145 ;
        RECT 394.185 56.765 394.565 57.145 ;
        RECT 404.470 56.765 404.850 57.145 ;
        RECT 414.760 56.765 415.140 57.145 ;
        RECT 425.045 56.765 425.425 57.145 ;
        RECT 426.465 56.765 426.845 57.145 ;
        RECT 436.755 56.765 437.135 57.145 ;
        RECT 447.040 56.765 447.420 57.145 ;
        RECT 457.330 56.765 457.710 57.145 ;
        RECT 467.615 56.765 467.995 57.145 ;
        RECT 469.035 56.765 469.415 57.145 ;
        RECT 479.325 56.765 479.705 57.145 ;
        RECT 489.610 56.765 489.990 57.145 ;
        RECT 499.900 56.765 500.280 57.145 ;
        RECT 510.185 56.765 510.565 57.145 ;
        RECT 511.605 56.765 511.985 57.145 ;
        RECT 521.895 56.765 522.275 57.145 ;
        RECT 532.180 56.765 532.560 57.145 ;
        RECT 542.470 56.765 542.850 57.145 ;
        RECT 552.755 56.765 553.135 57.145 ;
        RECT 554.175 56.765 554.555 57.145 ;
        RECT 564.465 56.765 564.845 57.145 ;
        RECT 574.750 56.765 575.130 57.145 ;
        RECT 585.040 56.765 585.420 57.145 ;
        RECT 595.325 56.765 595.705 57.145 ;
        RECT 596.745 56.765 597.125 57.145 ;
        RECT 607.035 56.765 607.415 57.145 ;
        RECT 617.320 56.765 617.700 57.145 ;
        RECT 627.610 56.765 627.990 57.145 ;
        RECT 637.895 56.765 638.275 57.145 ;
        RECT 639.315 56.765 639.695 57.145 ;
        RECT 649.605 56.765 649.985 57.145 ;
        RECT 659.890 56.765 660.270 57.145 ;
        RECT 670.180 56.765 670.560 57.145 ;
        RECT 680.465 56.765 680.845 57.145 ;
        RECT 0.765 56.105 1.145 56.485 ;
        RECT 11.055 56.105 11.435 56.485 ;
        RECT 21.340 56.105 21.720 56.485 ;
        RECT 31.630 56.105 32.010 56.485 ;
        RECT 41.915 56.105 42.295 56.485 ;
        RECT 43.335 56.105 43.715 56.485 ;
        RECT 53.625 56.105 54.005 56.485 ;
        RECT 63.910 56.105 64.290 56.485 ;
        RECT 74.200 56.105 74.580 56.485 ;
        RECT 84.485 56.105 84.865 56.485 ;
        RECT 85.905 56.105 86.285 56.485 ;
        RECT 96.195 56.105 96.575 56.485 ;
        RECT 106.480 56.105 106.860 56.485 ;
        RECT 116.770 56.105 117.150 56.485 ;
        RECT 127.055 56.105 127.435 56.485 ;
        RECT 128.475 56.105 128.855 56.485 ;
        RECT 138.765 56.105 139.145 56.485 ;
        RECT 149.050 56.105 149.430 56.485 ;
        RECT 159.340 56.105 159.720 56.485 ;
        RECT 169.625 56.105 170.005 56.485 ;
        RECT 171.045 56.105 171.425 56.485 ;
        RECT 181.335 56.105 181.715 56.485 ;
        RECT 191.620 56.105 192.000 56.485 ;
        RECT 201.910 56.105 202.290 56.485 ;
        RECT 212.195 56.105 212.575 56.485 ;
        RECT 213.615 56.105 213.995 56.485 ;
        RECT 223.905 56.105 224.285 56.485 ;
        RECT 234.190 56.105 234.570 56.485 ;
        RECT 244.480 56.105 244.860 56.485 ;
        RECT 254.765 56.105 255.145 56.485 ;
        RECT 256.185 56.105 256.565 56.485 ;
        RECT 266.475 56.105 266.855 56.485 ;
        RECT 276.760 56.105 277.140 56.485 ;
        RECT 287.050 56.105 287.430 56.485 ;
        RECT 297.335 56.105 297.715 56.485 ;
        RECT 298.755 56.105 299.135 56.485 ;
        RECT 309.045 56.105 309.425 56.485 ;
        RECT 319.330 56.105 319.710 56.485 ;
        RECT 329.620 56.105 330.000 56.485 ;
        RECT 339.905 56.105 340.285 56.485 ;
        RECT 341.325 56.105 341.705 56.485 ;
        RECT 351.615 56.105 351.995 56.485 ;
        RECT 361.900 56.105 362.280 56.485 ;
        RECT 372.190 56.105 372.570 56.485 ;
        RECT 382.475 56.105 382.855 56.485 ;
        RECT 383.895 56.105 384.275 56.485 ;
        RECT 394.185 56.105 394.565 56.485 ;
        RECT 404.470 56.105 404.850 56.485 ;
        RECT 414.760 56.105 415.140 56.485 ;
        RECT 425.045 56.105 425.425 56.485 ;
        RECT 426.465 56.105 426.845 56.485 ;
        RECT 436.755 56.105 437.135 56.485 ;
        RECT 447.040 56.105 447.420 56.485 ;
        RECT 457.330 56.105 457.710 56.485 ;
        RECT 467.615 56.105 467.995 56.485 ;
        RECT 469.035 56.105 469.415 56.485 ;
        RECT 479.325 56.105 479.705 56.485 ;
        RECT 489.610 56.105 489.990 56.485 ;
        RECT 499.900 56.105 500.280 56.485 ;
        RECT 510.185 56.105 510.565 56.485 ;
        RECT 511.605 56.105 511.985 56.485 ;
        RECT 521.895 56.105 522.275 56.485 ;
        RECT 532.180 56.105 532.560 56.485 ;
        RECT 542.470 56.105 542.850 56.485 ;
        RECT 552.755 56.105 553.135 56.485 ;
        RECT 554.175 56.105 554.555 56.485 ;
        RECT 564.465 56.105 564.845 56.485 ;
        RECT 574.750 56.105 575.130 56.485 ;
        RECT 585.040 56.105 585.420 56.485 ;
        RECT 595.325 56.105 595.705 56.485 ;
        RECT 596.745 56.105 597.125 56.485 ;
        RECT 607.035 56.105 607.415 56.485 ;
        RECT 617.320 56.105 617.700 56.485 ;
        RECT 627.610 56.105 627.990 56.485 ;
        RECT 637.895 56.105 638.275 56.485 ;
        RECT 639.315 56.105 639.695 56.485 ;
        RECT 649.605 56.105 649.985 56.485 ;
        RECT 659.890 56.105 660.270 56.485 ;
        RECT 670.180 56.105 670.560 56.485 ;
        RECT 680.465 56.105 680.845 56.485 ;
        RECT 0.765 55.445 1.145 55.825 ;
        RECT 11.055 55.445 11.435 55.825 ;
        RECT 21.340 55.445 21.720 55.825 ;
        RECT 31.630 55.445 32.010 55.825 ;
        RECT 41.915 55.445 42.295 55.825 ;
        RECT 43.335 55.445 43.715 55.825 ;
        RECT 53.625 55.445 54.005 55.825 ;
        RECT 63.910 55.445 64.290 55.825 ;
        RECT 74.200 55.445 74.580 55.825 ;
        RECT 84.485 55.445 84.865 55.825 ;
        RECT 85.905 55.445 86.285 55.825 ;
        RECT 96.195 55.445 96.575 55.825 ;
        RECT 106.480 55.445 106.860 55.825 ;
        RECT 116.770 55.445 117.150 55.825 ;
        RECT 127.055 55.445 127.435 55.825 ;
        RECT 128.475 55.445 128.855 55.825 ;
        RECT 138.765 55.445 139.145 55.825 ;
        RECT 149.050 55.445 149.430 55.825 ;
        RECT 159.340 55.445 159.720 55.825 ;
        RECT 169.625 55.445 170.005 55.825 ;
        RECT 171.045 55.445 171.425 55.825 ;
        RECT 181.335 55.445 181.715 55.825 ;
        RECT 191.620 55.445 192.000 55.825 ;
        RECT 201.910 55.445 202.290 55.825 ;
        RECT 212.195 55.445 212.575 55.825 ;
        RECT 213.615 55.445 213.995 55.825 ;
        RECT 223.905 55.445 224.285 55.825 ;
        RECT 234.190 55.445 234.570 55.825 ;
        RECT 244.480 55.445 244.860 55.825 ;
        RECT 254.765 55.445 255.145 55.825 ;
        RECT 256.185 55.445 256.565 55.825 ;
        RECT 266.475 55.445 266.855 55.825 ;
        RECT 276.760 55.445 277.140 55.825 ;
        RECT 287.050 55.445 287.430 55.825 ;
        RECT 297.335 55.445 297.715 55.825 ;
        RECT 298.755 55.445 299.135 55.825 ;
        RECT 309.045 55.445 309.425 55.825 ;
        RECT 319.330 55.445 319.710 55.825 ;
        RECT 329.620 55.445 330.000 55.825 ;
        RECT 339.905 55.445 340.285 55.825 ;
        RECT 341.325 55.445 341.705 55.825 ;
        RECT 351.615 55.445 351.995 55.825 ;
        RECT 361.900 55.445 362.280 55.825 ;
        RECT 372.190 55.445 372.570 55.825 ;
        RECT 382.475 55.445 382.855 55.825 ;
        RECT 383.895 55.445 384.275 55.825 ;
        RECT 394.185 55.445 394.565 55.825 ;
        RECT 404.470 55.445 404.850 55.825 ;
        RECT 414.760 55.445 415.140 55.825 ;
        RECT 425.045 55.445 425.425 55.825 ;
        RECT 426.465 55.445 426.845 55.825 ;
        RECT 436.755 55.445 437.135 55.825 ;
        RECT 447.040 55.445 447.420 55.825 ;
        RECT 457.330 55.445 457.710 55.825 ;
        RECT 467.615 55.445 467.995 55.825 ;
        RECT 469.035 55.445 469.415 55.825 ;
        RECT 479.325 55.445 479.705 55.825 ;
        RECT 489.610 55.445 489.990 55.825 ;
        RECT 499.900 55.445 500.280 55.825 ;
        RECT 510.185 55.445 510.565 55.825 ;
        RECT 511.605 55.445 511.985 55.825 ;
        RECT 521.895 55.445 522.275 55.825 ;
        RECT 532.180 55.445 532.560 55.825 ;
        RECT 542.470 55.445 542.850 55.825 ;
        RECT 552.755 55.445 553.135 55.825 ;
        RECT 554.175 55.445 554.555 55.825 ;
        RECT 564.465 55.445 564.845 55.825 ;
        RECT 574.750 55.445 575.130 55.825 ;
        RECT 585.040 55.445 585.420 55.825 ;
        RECT 595.325 55.445 595.705 55.825 ;
        RECT 596.745 55.445 597.125 55.825 ;
        RECT 607.035 55.445 607.415 55.825 ;
        RECT 617.320 55.445 617.700 55.825 ;
        RECT 627.610 55.445 627.990 55.825 ;
        RECT 637.895 55.445 638.275 55.825 ;
        RECT 639.315 55.445 639.695 55.825 ;
        RECT 649.605 55.445 649.985 55.825 ;
        RECT 659.890 55.445 660.270 55.825 ;
        RECT 670.180 55.445 670.560 55.825 ;
        RECT 680.465 55.445 680.845 55.825 ;
        RECT 0.765 54.785 1.145 55.165 ;
        RECT 11.055 54.785 11.435 55.165 ;
        RECT 21.340 54.785 21.720 55.165 ;
        RECT 31.630 54.785 32.010 55.165 ;
        RECT 41.915 54.785 42.295 55.165 ;
        RECT 43.335 54.785 43.715 55.165 ;
        RECT 53.625 54.785 54.005 55.165 ;
        RECT 63.910 54.785 64.290 55.165 ;
        RECT 74.200 54.785 74.580 55.165 ;
        RECT 84.485 54.785 84.865 55.165 ;
        RECT 85.905 54.785 86.285 55.165 ;
        RECT 96.195 54.785 96.575 55.165 ;
        RECT 106.480 54.785 106.860 55.165 ;
        RECT 116.770 54.785 117.150 55.165 ;
        RECT 127.055 54.785 127.435 55.165 ;
        RECT 128.475 54.785 128.855 55.165 ;
        RECT 138.765 54.785 139.145 55.165 ;
        RECT 149.050 54.785 149.430 55.165 ;
        RECT 159.340 54.785 159.720 55.165 ;
        RECT 169.625 54.785 170.005 55.165 ;
        RECT 171.045 54.785 171.425 55.165 ;
        RECT 181.335 54.785 181.715 55.165 ;
        RECT 191.620 54.785 192.000 55.165 ;
        RECT 201.910 54.785 202.290 55.165 ;
        RECT 212.195 54.785 212.575 55.165 ;
        RECT 213.615 54.785 213.995 55.165 ;
        RECT 223.905 54.785 224.285 55.165 ;
        RECT 234.190 54.785 234.570 55.165 ;
        RECT 244.480 54.785 244.860 55.165 ;
        RECT 254.765 54.785 255.145 55.165 ;
        RECT 256.185 54.785 256.565 55.165 ;
        RECT 266.475 54.785 266.855 55.165 ;
        RECT 276.760 54.785 277.140 55.165 ;
        RECT 287.050 54.785 287.430 55.165 ;
        RECT 297.335 54.785 297.715 55.165 ;
        RECT 298.755 54.785 299.135 55.165 ;
        RECT 309.045 54.785 309.425 55.165 ;
        RECT 319.330 54.785 319.710 55.165 ;
        RECT 329.620 54.785 330.000 55.165 ;
        RECT 339.905 54.785 340.285 55.165 ;
        RECT 341.325 54.785 341.705 55.165 ;
        RECT 351.615 54.785 351.995 55.165 ;
        RECT 361.900 54.785 362.280 55.165 ;
        RECT 372.190 54.785 372.570 55.165 ;
        RECT 382.475 54.785 382.855 55.165 ;
        RECT 383.895 54.785 384.275 55.165 ;
        RECT 394.185 54.785 394.565 55.165 ;
        RECT 404.470 54.785 404.850 55.165 ;
        RECT 414.760 54.785 415.140 55.165 ;
        RECT 425.045 54.785 425.425 55.165 ;
        RECT 426.465 54.785 426.845 55.165 ;
        RECT 436.755 54.785 437.135 55.165 ;
        RECT 447.040 54.785 447.420 55.165 ;
        RECT 457.330 54.785 457.710 55.165 ;
        RECT 467.615 54.785 467.995 55.165 ;
        RECT 469.035 54.785 469.415 55.165 ;
        RECT 479.325 54.785 479.705 55.165 ;
        RECT 489.610 54.785 489.990 55.165 ;
        RECT 499.900 54.785 500.280 55.165 ;
        RECT 510.185 54.785 510.565 55.165 ;
        RECT 511.605 54.785 511.985 55.165 ;
        RECT 521.895 54.785 522.275 55.165 ;
        RECT 532.180 54.785 532.560 55.165 ;
        RECT 542.470 54.785 542.850 55.165 ;
        RECT 552.755 54.785 553.135 55.165 ;
        RECT 554.175 54.785 554.555 55.165 ;
        RECT 564.465 54.785 564.845 55.165 ;
        RECT 574.750 54.785 575.130 55.165 ;
        RECT 585.040 54.785 585.420 55.165 ;
        RECT 595.325 54.785 595.705 55.165 ;
        RECT 596.745 54.785 597.125 55.165 ;
        RECT 607.035 54.785 607.415 55.165 ;
        RECT 617.320 54.785 617.700 55.165 ;
        RECT 627.610 54.785 627.990 55.165 ;
        RECT 637.895 54.785 638.275 55.165 ;
        RECT 639.315 54.785 639.695 55.165 ;
        RECT 649.605 54.785 649.985 55.165 ;
        RECT 659.890 54.785 660.270 55.165 ;
        RECT 670.180 54.785 670.560 55.165 ;
        RECT 680.465 54.785 680.845 55.165 ;
        RECT 682.310 55.115 682.690 55.495 ;
        RECT 684.095 55.115 684.475 55.495 ;
        RECT 686.950 55.115 687.330 55.495 ;
        RECT 688.735 55.115 689.115 55.495 ;
        RECT 691.590 55.115 691.970 55.495 ;
        RECT 693.375 55.115 693.755 55.495 ;
        RECT 696.230 55.115 696.610 55.495 ;
        RECT 698.015 55.115 698.395 55.495 ;
        RECT 700.870 55.115 701.250 55.495 ;
        RECT 702.655 55.115 703.035 55.495 ;
        RECT 705.510 55.115 705.890 55.495 ;
        RECT 707.295 55.115 707.675 55.495 ;
        RECT 710.150 55.115 710.530 55.495 ;
        RECT 711.935 55.115 712.315 55.495 ;
        RECT 714.790 55.115 715.170 55.495 ;
        RECT 716.575 55.115 716.955 55.495 ;
        RECT 0.765 54.125 1.145 54.505 ;
        RECT 11.055 54.125 11.435 54.505 ;
        RECT 21.340 54.125 21.720 54.505 ;
        RECT 31.630 54.125 32.010 54.505 ;
        RECT 41.915 54.125 42.295 54.505 ;
        RECT 43.335 54.125 43.715 54.505 ;
        RECT 53.625 54.125 54.005 54.505 ;
        RECT 63.910 54.125 64.290 54.505 ;
        RECT 74.200 54.125 74.580 54.505 ;
        RECT 84.485 54.125 84.865 54.505 ;
        RECT 85.905 54.125 86.285 54.505 ;
        RECT 96.195 54.125 96.575 54.505 ;
        RECT 106.480 54.125 106.860 54.505 ;
        RECT 116.770 54.125 117.150 54.505 ;
        RECT 127.055 54.125 127.435 54.505 ;
        RECT 128.475 54.125 128.855 54.505 ;
        RECT 138.765 54.125 139.145 54.505 ;
        RECT 149.050 54.125 149.430 54.505 ;
        RECT 159.340 54.125 159.720 54.505 ;
        RECT 169.625 54.125 170.005 54.505 ;
        RECT 171.045 54.125 171.425 54.505 ;
        RECT 181.335 54.125 181.715 54.505 ;
        RECT 191.620 54.125 192.000 54.505 ;
        RECT 201.910 54.125 202.290 54.505 ;
        RECT 212.195 54.125 212.575 54.505 ;
        RECT 213.615 54.125 213.995 54.505 ;
        RECT 223.905 54.125 224.285 54.505 ;
        RECT 234.190 54.125 234.570 54.505 ;
        RECT 244.480 54.125 244.860 54.505 ;
        RECT 254.765 54.125 255.145 54.505 ;
        RECT 256.185 54.125 256.565 54.505 ;
        RECT 266.475 54.125 266.855 54.505 ;
        RECT 276.760 54.125 277.140 54.505 ;
        RECT 287.050 54.125 287.430 54.505 ;
        RECT 297.335 54.125 297.715 54.505 ;
        RECT 298.755 54.125 299.135 54.505 ;
        RECT 309.045 54.125 309.425 54.505 ;
        RECT 319.330 54.125 319.710 54.505 ;
        RECT 329.620 54.125 330.000 54.505 ;
        RECT 339.905 54.125 340.285 54.505 ;
        RECT 341.325 54.125 341.705 54.505 ;
        RECT 351.615 54.125 351.995 54.505 ;
        RECT 361.900 54.125 362.280 54.505 ;
        RECT 372.190 54.125 372.570 54.505 ;
        RECT 382.475 54.125 382.855 54.505 ;
        RECT 383.895 54.125 384.275 54.505 ;
        RECT 394.185 54.125 394.565 54.505 ;
        RECT 404.470 54.125 404.850 54.505 ;
        RECT 414.760 54.125 415.140 54.505 ;
        RECT 425.045 54.125 425.425 54.505 ;
        RECT 426.465 54.125 426.845 54.505 ;
        RECT 436.755 54.125 437.135 54.505 ;
        RECT 447.040 54.125 447.420 54.505 ;
        RECT 457.330 54.125 457.710 54.505 ;
        RECT 467.615 54.125 467.995 54.505 ;
        RECT 469.035 54.125 469.415 54.505 ;
        RECT 479.325 54.125 479.705 54.505 ;
        RECT 489.610 54.125 489.990 54.505 ;
        RECT 499.900 54.125 500.280 54.505 ;
        RECT 510.185 54.125 510.565 54.505 ;
        RECT 511.605 54.125 511.985 54.505 ;
        RECT 521.895 54.125 522.275 54.505 ;
        RECT 532.180 54.125 532.560 54.505 ;
        RECT 542.470 54.125 542.850 54.505 ;
        RECT 552.755 54.125 553.135 54.505 ;
        RECT 554.175 54.125 554.555 54.505 ;
        RECT 564.465 54.125 564.845 54.505 ;
        RECT 574.750 54.125 575.130 54.505 ;
        RECT 585.040 54.125 585.420 54.505 ;
        RECT 595.325 54.125 595.705 54.505 ;
        RECT 596.745 54.125 597.125 54.505 ;
        RECT 607.035 54.125 607.415 54.505 ;
        RECT 617.320 54.125 617.700 54.505 ;
        RECT 627.610 54.125 627.990 54.505 ;
        RECT 637.895 54.125 638.275 54.505 ;
        RECT 639.315 54.125 639.695 54.505 ;
        RECT 649.605 54.125 649.985 54.505 ;
        RECT 659.890 54.125 660.270 54.505 ;
        RECT 670.180 54.125 670.560 54.505 ;
        RECT 680.465 54.125 680.845 54.505 ;
        RECT 682.310 54.455 682.690 54.835 ;
        RECT 684.095 54.455 684.475 54.835 ;
        RECT 686.950 54.455 687.330 54.835 ;
        RECT 688.735 54.455 689.115 54.835 ;
        RECT 691.590 54.455 691.970 54.835 ;
        RECT 693.375 54.455 693.755 54.835 ;
        RECT 696.230 54.455 696.610 54.835 ;
        RECT 698.015 54.455 698.395 54.835 ;
        RECT 700.870 54.455 701.250 54.835 ;
        RECT 702.655 54.455 703.035 54.835 ;
        RECT 705.510 54.455 705.890 54.835 ;
        RECT 707.295 54.455 707.675 54.835 ;
        RECT 710.150 54.455 710.530 54.835 ;
        RECT 711.935 54.455 712.315 54.835 ;
        RECT 714.790 54.455 715.170 54.835 ;
        RECT 716.575 54.455 716.955 54.835 ;
        RECT 0.765 53.465 1.145 53.845 ;
        RECT 11.055 53.465 11.435 53.845 ;
        RECT 21.340 53.465 21.720 53.845 ;
        RECT 31.630 53.465 32.010 53.845 ;
        RECT 41.915 53.465 42.295 53.845 ;
        RECT 43.335 53.465 43.715 53.845 ;
        RECT 53.625 53.465 54.005 53.845 ;
        RECT 63.910 53.465 64.290 53.845 ;
        RECT 74.200 53.465 74.580 53.845 ;
        RECT 84.485 53.465 84.865 53.845 ;
        RECT 85.905 53.465 86.285 53.845 ;
        RECT 96.195 53.465 96.575 53.845 ;
        RECT 106.480 53.465 106.860 53.845 ;
        RECT 116.770 53.465 117.150 53.845 ;
        RECT 127.055 53.465 127.435 53.845 ;
        RECT 128.475 53.465 128.855 53.845 ;
        RECT 138.765 53.465 139.145 53.845 ;
        RECT 149.050 53.465 149.430 53.845 ;
        RECT 159.340 53.465 159.720 53.845 ;
        RECT 169.625 53.465 170.005 53.845 ;
        RECT 171.045 53.465 171.425 53.845 ;
        RECT 181.335 53.465 181.715 53.845 ;
        RECT 191.620 53.465 192.000 53.845 ;
        RECT 201.910 53.465 202.290 53.845 ;
        RECT 212.195 53.465 212.575 53.845 ;
        RECT 213.615 53.465 213.995 53.845 ;
        RECT 223.905 53.465 224.285 53.845 ;
        RECT 234.190 53.465 234.570 53.845 ;
        RECT 244.480 53.465 244.860 53.845 ;
        RECT 254.765 53.465 255.145 53.845 ;
        RECT 256.185 53.465 256.565 53.845 ;
        RECT 266.475 53.465 266.855 53.845 ;
        RECT 276.760 53.465 277.140 53.845 ;
        RECT 287.050 53.465 287.430 53.845 ;
        RECT 297.335 53.465 297.715 53.845 ;
        RECT 298.755 53.465 299.135 53.845 ;
        RECT 309.045 53.465 309.425 53.845 ;
        RECT 319.330 53.465 319.710 53.845 ;
        RECT 329.620 53.465 330.000 53.845 ;
        RECT 339.905 53.465 340.285 53.845 ;
        RECT 341.325 53.465 341.705 53.845 ;
        RECT 351.615 53.465 351.995 53.845 ;
        RECT 361.900 53.465 362.280 53.845 ;
        RECT 372.190 53.465 372.570 53.845 ;
        RECT 382.475 53.465 382.855 53.845 ;
        RECT 383.895 53.465 384.275 53.845 ;
        RECT 394.185 53.465 394.565 53.845 ;
        RECT 404.470 53.465 404.850 53.845 ;
        RECT 414.760 53.465 415.140 53.845 ;
        RECT 425.045 53.465 425.425 53.845 ;
        RECT 426.465 53.465 426.845 53.845 ;
        RECT 436.755 53.465 437.135 53.845 ;
        RECT 447.040 53.465 447.420 53.845 ;
        RECT 457.330 53.465 457.710 53.845 ;
        RECT 467.615 53.465 467.995 53.845 ;
        RECT 469.035 53.465 469.415 53.845 ;
        RECT 479.325 53.465 479.705 53.845 ;
        RECT 489.610 53.465 489.990 53.845 ;
        RECT 499.900 53.465 500.280 53.845 ;
        RECT 510.185 53.465 510.565 53.845 ;
        RECT 511.605 53.465 511.985 53.845 ;
        RECT 521.895 53.465 522.275 53.845 ;
        RECT 532.180 53.465 532.560 53.845 ;
        RECT 542.470 53.465 542.850 53.845 ;
        RECT 552.755 53.465 553.135 53.845 ;
        RECT 554.175 53.465 554.555 53.845 ;
        RECT 564.465 53.465 564.845 53.845 ;
        RECT 574.750 53.465 575.130 53.845 ;
        RECT 585.040 53.465 585.420 53.845 ;
        RECT 595.325 53.465 595.705 53.845 ;
        RECT 596.745 53.465 597.125 53.845 ;
        RECT 607.035 53.465 607.415 53.845 ;
        RECT 617.320 53.465 617.700 53.845 ;
        RECT 627.610 53.465 627.990 53.845 ;
        RECT 637.895 53.465 638.275 53.845 ;
        RECT 639.315 53.465 639.695 53.845 ;
        RECT 649.605 53.465 649.985 53.845 ;
        RECT 659.890 53.465 660.270 53.845 ;
        RECT 670.180 53.465 670.560 53.845 ;
        RECT 680.465 53.465 680.845 53.845 ;
        RECT 682.310 53.795 682.690 54.175 ;
        RECT 684.095 53.795 684.475 54.175 ;
        RECT 686.950 53.795 687.330 54.175 ;
        RECT 688.735 53.795 689.115 54.175 ;
        RECT 691.590 53.795 691.970 54.175 ;
        RECT 693.375 53.795 693.755 54.175 ;
        RECT 696.230 53.795 696.610 54.175 ;
        RECT 698.015 53.795 698.395 54.175 ;
        RECT 700.870 53.795 701.250 54.175 ;
        RECT 702.655 53.795 703.035 54.175 ;
        RECT 705.510 53.795 705.890 54.175 ;
        RECT 707.295 53.795 707.675 54.175 ;
        RECT 710.150 53.795 710.530 54.175 ;
        RECT 711.935 53.795 712.315 54.175 ;
        RECT 714.790 53.795 715.170 54.175 ;
        RECT 716.575 53.795 716.955 54.175 ;
        RECT 0.765 52.805 1.145 53.185 ;
        RECT 11.055 52.805 11.435 53.185 ;
        RECT 21.340 52.805 21.720 53.185 ;
        RECT 31.630 52.805 32.010 53.185 ;
        RECT 41.915 52.805 42.295 53.185 ;
        RECT 43.335 52.805 43.715 53.185 ;
        RECT 53.625 52.805 54.005 53.185 ;
        RECT 63.910 52.805 64.290 53.185 ;
        RECT 74.200 52.805 74.580 53.185 ;
        RECT 84.485 52.805 84.865 53.185 ;
        RECT 85.905 52.805 86.285 53.185 ;
        RECT 96.195 52.805 96.575 53.185 ;
        RECT 106.480 52.805 106.860 53.185 ;
        RECT 116.770 52.805 117.150 53.185 ;
        RECT 127.055 52.805 127.435 53.185 ;
        RECT 128.475 52.805 128.855 53.185 ;
        RECT 138.765 52.805 139.145 53.185 ;
        RECT 149.050 52.805 149.430 53.185 ;
        RECT 159.340 52.805 159.720 53.185 ;
        RECT 169.625 52.805 170.005 53.185 ;
        RECT 171.045 52.805 171.425 53.185 ;
        RECT 181.335 52.805 181.715 53.185 ;
        RECT 191.620 52.805 192.000 53.185 ;
        RECT 201.910 52.805 202.290 53.185 ;
        RECT 212.195 52.805 212.575 53.185 ;
        RECT 213.615 52.805 213.995 53.185 ;
        RECT 223.905 52.805 224.285 53.185 ;
        RECT 234.190 52.805 234.570 53.185 ;
        RECT 244.480 52.805 244.860 53.185 ;
        RECT 254.765 52.805 255.145 53.185 ;
        RECT 256.185 52.805 256.565 53.185 ;
        RECT 266.475 52.805 266.855 53.185 ;
        RECT 276.760 52.805 277.140 53.185 ;
        RECT 287.050 52.805 287.430 53.185 ;
        RECT 297.335 52.805 297.715 53.185 ;
        RECT 298.755 52.805 299.135 53.185 ;
        RECT 309.045 52.805 309.425 53.185 ;
        RECT 319.330 52.805 319.710 53.185 ;
        RECT 329.620 52.805 330.000 53.185 ;
        RECT 339.905 52.805 340.285 53.185 ;
        RECT 341.325 52.805 341.705 53.185 ;
        RECT 351.615 52.805 351.995 53.185 ;
        RECT 361.900 52.805 362.280 53.185 ;
        RECT 372.190 52.805 372.570 53.185 ;
        RECT 382.475 52.805 382.855 53.185 ;
        RECT 383.895 52.805 384.275 53.185 ;
        RECT 394.185 52.805 394.565 53.185 ;
        RECT 404.470 52.805 404.850 53.185 ;
        RECT 414.760 52.805 415.140 53.185 ;
        RECT 425.045 52.805 425.425 53.185 ;
        RECT 426.465 52.805 426.845 53.185 ;
        RECT 436.755 52.805 437.135 53.185 ;
        RECT 447.040 52.805 447.420 53.185 ;
        RECT 457.330 52.805 457.710 53.185 ;
        RECT 467.615 52.805 467.995 53.185 ;
        RECT 469.035 52.805 469.415 53.185 ;
        RECT 479.325 52.805 479.705 53.185 ;
        RECT 489.610 52.805 489.990 53.185 ;
        RECT 499.900 52.805 500.280 53.185 ;
        RECT 510.185 52.805 510.565 53.185 ;
        RECT 511.605 52.805 511.985 53.185 ;
        RECT 521.895 52.805 522.275 53.185 ;
        RECT 532.180 52.805 532.560 53.185 ;
        RECT 542.470 52.805 542.850 53.185 ;
        RECT 552.755 52.805 553.135 53.185 ;
        RECT 554.175 52.805 554.555 53.185 ;
        RECT 564.465 52.805 564.845 53.185 ;
        RECT 574.750 52.805 575.130 53.185 ;
        RECT 585.040 52.805 585.420 53.185 ;
        RECT 595.325 52.805 595.705 53.185 ;
        RECT 596.745 52.805 597.125 53.185 ;
        RECT 607.035 52.805 607.415 53.185 ;
        RECT 617.320 52.805 617.700 53.185 ;
        RECT 627.610 52.805 627.990 53.185 ;
        RECT 637.895 52.805 638.275 53.185 ;
        RECT 639.315 52.805 639.695 53.185 ;
        RECT 649.605 52.805 649.985 53.185 ;
        RECT 659.890 52.805 660.270 53.185 ;
        RECT 670.180 52.805 670.560 53.185 ;
        RECT 680.465 52.805 680.845 53.185 ;
        RECT 682.310 53.135 682.690 53.515 ;
        RECT 684.095 53.135 684.475 53.515 ;
        RECT 686.950 53.135 687.330 53.515 ;
        RECT 688.735 53.135 689.115 53.515 ;
        RECT 691.590 53.135 691.970 53.515 ;
        RECT 693.375 53.135 693.755 53.515 ;
        RECT 696.230 53.135 696.610 53.515 ;
        RECT 698.015 53.135 698.395 53.515 ;
        RECT 700.870 53.135 701.250 53.515 ;
        RECT 702.655 53.135 703.035 53.515 ;
        RECT 705.510 53.135 705.890 53.515 ;
        RECT 707.295 53.135 707.675 53.515 ;
        RECT 710.150 53.135 710.530 53.515 ;
        RECT 711.935 53.135 712.315 53.515 ;
        RECT 714.790 53.135 715.170 53.515 ;
        RECT 716.575 53.135 716.955 53.515 ;
        RECT 0.765 52.145 1.145 52.525 ;
        RECT 11.055 52.145 11.435 52.525 ;
        RECT 21.340 52.145 21.720 52.525 ;
        RECT 31.630 52.145 32.010 52.525 ;
        RECT 41.915 52.145 42.295 52.525 ;
        RECT 43.335 52.145 43.715 52.525 ;
        RECT 53.625 52.145 54.005 52.525 ;
        RECT 63.910 52.145 64.290 52.525 ;
        RECT 74.200 52.145 74.580 52.525 ;
        RECT 84.485 52.145 84.865 52.525 ;
        RECT 85.905 52.145 86.285 52.525 ;
        RECT 96.195 52.145 96.575 52.525 ;
        RECT 106.480 52.145 106.860 52.525 ;
        RECT 116.770 52.145 117.150 52.525 ;
        RECT 127.055 52.145 127.435 52.525 ;
        RECT 128.475 52.145 128.855 52.525 ;
        RECT 138.765 52.145 139.145 52.525 ;
        RECT 149.050 52.145 149.430 52.525 ;
        RECT 159.340 52.145 159.720 52.525 ;
        RECT 169.625 52.145 170.005 52.525 ;
        RECT 171.045 52.145 171.425 52.525 ;
        RECT 181.335 52.145 181.715 52.525 ;
        RECT 191.620 52.145 192.000 52.525 ;
        RECT 201.910 52.145 202.290 52.525 ;
        RECT 212.195 52.145 212.575 52.525 ;
        RECT 213.615 52.145 213.995 52.525 ;
        RECT 223.905 52.145 224.285 52.525 ;
        RECT 234.190 52.145 234.570 52.525 ;
        RECT 244.480 52.145 244.860 52.525 ;
        RECT 254.765 52.145 255.145 52.525 ;
        RECT 256.185 52.145 256.565 52.525 ;
        RECT 266.475 52.145 266.855 52.525 ;
        RECT 276.760 52.145 277.140 52.525 ;
        RECT 287.050 52.145 287.430 52.525 ;
        RECT 297.335 52.145 297.715 52.525 ;
        RECT 298.755 52.145 299.135 52.525 ;
        RECT 309.045 52.145 309.425 52.525 ;
        RECT 319.330 52.145 319.710 52.525 ;
        RECT 329.620 52.145 330.000 52.525 ;
        RECT 339.905 52.145 340.285 52.525 ;
        RECT 341.325 52.145 341.705 52.525 ;
        RECT 351.615 52.145 351.995 52.525 ;
        RECT 361.900 52.145 362.280 52.525 ;
        RECT 372.190 52.145 372.570 52.525 ;
        RECT 382.475 52.145 382.855 52.525 ;
        RECT 383.895 52.145 384.275 52.525 ;
        RECT 394.185 52.145 394.565 52.525 ;
        RECT 404.470 52.145 404.850 52.525 ;
        RECT 414.760 52.145 415.140 52.525 ;
        RECT 425.045 52.145 425.425 52.525 ;
        RECT 426.465 52.145 426.845 52.525 ;
        RECT 436.755 52.145 437.135 52.525 ;
        RECT 447.040 52.145 447.420 52.525 ;
        RECT 457.330 52.145 457.710 52.525 ;
        RECT 467.615 52.145 467.995 52.525 ;
        RECT 469.035 52.145 469.415 52.525 ;
        RECT 479.325 52.145 479.705 52.525 ;
        RECT 489.610 52.145 489.990 52.525 ;
        RECT 499.900 52.145 500.280 52.525 ;
        RECT 510.185 52.145 510.565 52.525 ;
        RECT 511.605 52.145 511.985 52.525 ;
        RECT 521.895 52.145 522.275 52.525 ;
        RECT 532.180 52.145 532.560 52.525 ;
        RECT 542.470 52.145 542.850 52.525 ;
        RECT 552.755 52.145 553.135 52.525 ;
        RECT 554.175 52.145 554.555 52.525 ;
        RECT 564.465 52.145 564.845 52.525 ;
        RECT 574.750 52.145 575.130 52.525 ;
        RECT 585.040 52.145 585.420 52.525 ;
        RECT 595.325 52.145 595.705 52.525 ;
        RECT 596.745 52.145 597.125 52.525 ;
        RECT 607.035 52.145 607.415 52.525 ;
        RECT 617.320 52.145 617.700 52.525 ;
        RECT 627.610 52.145 627.990 52.525 ;
        RECT 637.895 52.145 638.275 52.525 ;
        RECT 639.315 52.145 639.695 52.525 ;
        RECT 649.605 52.145 649.985 52.525 ;
        RECT 659.890 52.145 660.270 52.525 ;
        RECT 670.180 52.145 670.560 52.525 ;
        RECT 680.465 52.145 680.845 52.525 ;
        RECT 682.310 52.475 682.690 52.855 ;
        RECT 684.095 52.475 684.475 52.855 ;
        RECT 686.950 52.475 687.330 52.855 ;
        RECT 688.735 52.475 689.115 52.855 ;
        RECT 691.590 52.475 691.970 52.855 ;
        RECT 693.375 52.475 693.755 52.855 ;
        RECT 696.230 52.475 696.610 52.855 ;
        RECT 698.015 52.475 698.395 52.855 ;
        RECT 700.870 52.475 701.250 52.855 ;
        RECT 702.655 52.475 703.035 52.855 ;
        RECT 705.510 52.475 705.890 52.855 ;
        RECT 707.295 52.475 707.675 52.855 ;
        RECT 710.150 52.475 710.530 52.855 ;
        RECT 711.935 52.475 712.315 52.855 ;
        RECT 714.790 52.475 715.170 52.855 ;
        RECT 716.575 52.475 716.955 52.855 ;
        RECT 0.765 51.485 1.145 51.865 ;
        RECT 11.055 51.485 11.435 51.865 ;
        RECT 21.340 51.485 21.720 51.865 ;
        RECT 31.630 51.485 32.010 51.865 ;
        RECT 41.915 51.485 42.295 51.865 ;
        RECT 43.335 51.485 43.715 51.865 ;
        RECT 53.625 51.485 54.005 51.865 ;
        RECT 63.910 51.485 64.290 51.865 ;
        RECT 74.200 51.485 74.580 51.865 ;
        RECT 84.485 51.485 84.865 51.865 ;
        RECT 85.905 51.485 86.285 51.865 ;
        RECT 96.195 51.485 96.575 51.865 ;
        RECT 106.480 51.485 106.860 51.865 ;
        RECT 116.770 51.485 117.150 51.865 ;
        RECT 127.055 51.485 127.435 51.865 ;
        RECT 128.475 51.485 128.855 51.865 ;
        RECT 138.765 51.485 139.145 51.865 ;
        RECT 149.050 51.485 149.430 51.865 ;
        RECT 159.340 51.485 159.720 51.865 ;
        RECT 169.625 51.485 170.005 51.865 ;
        RECT 171.045 51.485 171.425 51.865 ;
        RECT 181.335 51.485 181.715 51.865 ;
        RECT 191.620 51.485 192.000 51.865 ;
        RECT 201.910 51.485 202.290 51.865 ;
        RECT 212.195 51.485 212.575 51.865 ;
        RECT 213.615 51.485 213.995 51.865 ;
        RECT 223.905 51.485 224.285 51.865 ;
        RECT 234.190 51.485 234.570 51.865 ;
        RECT 244.480 51.485 244.860 51.865 ;
        RECT 254.765 51.485 255.145 51.865 ;
        RECT 256.185 51.485 256.565 51.865 ;
        RECT 266.475 51.485 266.855 51.865 ;
        RECT 276.760 51.485 277.140 51.865 ;
        RECT 287.050 51.485 287.430 51.865 ;
        RECT 297.335 51.485 297.715 51.865 ;
        RECT 298.755 51.485 299.135 51.865 ;
        RECT 309.045 51.485 309.425 51.865 ;
        RECT 319.330 51.485 319.710 51.865 ;
        RECT 329.620 51.485 330.000 51.865 ;
        RECT 339.905 51.485 340.285 51.865 ;
        RECT 341.325 51.485 341.705 51.865 ;
        RECT 351.615 51.485 351.995 51.865 ;
        RECT 361.900 51.485 362.280 51.865 ;
        RECT 372.190 51.485 372.570 51.865 ;
        RECT 382.475 51.485 382.855 51.865 ;
        RECT 383.895 51.485 384.275 51.865 ;
        RECT 394.185 51.485 394.565 51.865 ;
        RECT 404.470 51.485 404.850 51.865 ;
        RECT 414.760 51.485 415.140 51.865 ;
        RECT 425.045 51.485 425.425 51.865 ;
        RECT 426.465 51.485 426.845 51.865 ;
        RECT 436.755 51.485 437.135 51.865 ;
        RECT 447.040 51.485 447.420 51.865 ;
        RECT 457.330 51.485 457.710 51.865 ;
        RECT 467.615 51.485 467.995 51.865 ;
        RECT 469.035 51.485 469.415 51.865 ;
        RECT 479.325 51.485 479.705 51.865 ;
        RECT 489.610 51.485 489.990 51.865 ;
        RECT 499.900 51.485 500.280 51.865 ;
        RECT 510.185 51.485 510.565 51.865 ;
        RECT 511.605 51.485 511.985 51.865 ;
        RECT 521.895 51.485 522.275 51.865 ;
        RECT 532.180 51.485 532.560 51.865 ;
        RECT 542.470 51.485 542.850 51.865 ;
        RECT 552.755 51.485 553.135 51.865 ;
        RECT 554.175 51.485 554.555 51.865 ;
        RECT 564.465 51.485 564.845 51.865 ;
        RECT 574.750 51.485 575.130 51.865 ;
        RECT 585.040 51.485 585.420 51.865 ;
        RECT 595.325 51.485 595.705 51.865 ;
        RECT 596.745 51.485 597.125 51.865 ;
        RECT 607.035 51.485 607.415 51.865 ;
        RECT 617.320 51.485 617.700 51.865 ;
        RECT 627.610 51.485 627.990 51.865 ;
        RECT 637.895 51.485 638.275 51.865 ;
        RECT 639.315 51.485 639.695 51.865 ;
        RECT 649.605 51.485 649.985 51.865 ;
        RECT 659.890 51.485 660.270 51.865 ;
        RECT 670.180 51.485 670.560 51.865 ;
        RECT 680.465 51.485 680.845 51.865 ;
        RECT 682.310 51.815 682.690 52.195 ;
        RECT 684.095 51.815 684.475 52.195 ;
        RECT 686.950 51.815 687.330 52.195 ;
        RECT 688.735 51.815 689.115 52.195 ;
        RECT 691.590 51.815 691.970 52.195 ;
        RECT 693.375 51.815 693.755 52.195 ;
        RECT 696.230 51.815 696.610 52.195 ;
        RECT 698.015 51.815 698.395 52.195 ;
        RECT 700.870 51.815 701.250 52.195 ;
        RECT 702.655 51.815 703.035 52.195 ;
        RECT 705.510 51.815 705.890 52.195 ;
        RECT 707.295 51.815 707.675 52.195 ;
        RECT 710.150 51.815 710.530 52.195 ;
        RECT 711.935 51.815 712.315 52.195 ;
        RECT 714.790 51.815 715.170 52.195 ;
        RECT 716.575 51.815 716.955 52.195 ;
        RECT 0.765 50.825 1.145 51.205 ;
        RECT 11.055 50.825 11.435 51.205 ;
        RECT 21.340 50.825 21.720 51.205 ;
        RECT 31.630 50.825 32.010 51.205 ;
        RECT 41.915 50.825 42.295 51.205 ;
        RECT 43.335 50.825 43.715 51.205 ;
        RECT 53.625 50.825 54.005 51.205 ;
        RECT 63.910 50.825 64.290 51.205 ;
        RECT 74.200 50.825 74.580 51.205 ;
        RECT 84.485 50.825 84.865 51.205 ;
        RECT 85.905 50.825 86.285 51.205 ;
        RECT 96.195 50.825 96.575 51.205 ;
        RECT 106.480 50.825 106.860 51.205 ;
        RECT 116.770 50.825 117.150 51.205 ;
        RECT 127.055 50.825 127.435 51.205 ;
        RECT 128.475 50.825 128.855 51.205 ;
        RECT 138.765 50.825 139.145 51.205 ;
        RECT 149.050 50.825 149.430 51.205 ;
        RECT 159.340 50.825 159.720 51.205 ;
        RECT 169.625 50.825 170.005 51.205 ;
        RECT 171.045 50.825 171.425 51.205 ;
        RECT 181.335 50.825 181.715 51.205 ;
        RECT 191.620 50.825 192.000 51.205 ;
        RECT 201.910 50.825 202.290 51.205 ;
        RECT 212.195 50.825 212.575 51.205 ;
        RECT 213.615 50.825 213.995 51.205 ;
        RECT 223.905 50.825 224.285 51.205 ;
        RECT 234.190 50.825 234.570 51.205 ;
        RECT 244.480 50.825 244.860 51.205 ;
        RECT 254.765 50.825 255.145 51.205 ;
        RECT 256.185 50.825 256.565 51.205 ;
        RECT 266.475 50.825 266.855 51.205 ;
        RECT 276.760 50.825 277.140 51.205 ;
        RECT 287.050 50.825 287.430 51.205 ;
        RECT 297.335 50.825 297.715 51.205 ;
        RECT 298.755 50.825 299.135 51.205 ;
        RECT 309.045 50.825 309.425 51.205 ;
        RECT 319.330 50.825 319.710 51.205 ;
        RECT 329.620 50.825 330.000 51.205 ;
        RECT 339.905 50.825 340.285 51.205 ;
        RECT 341.325 50.825 341.705 51.205 ;
        RECT 351.615 50.825 351.995 51.205 ;
        RECT 361.900 50.825 362.280 51.205 ;
        RECT 372.190 50.825 372.570 51.205 ;
        RECT 382.475 50.825 382.855 51.205 ;
        RECT 383.895 50.825 384.275 51.205 ;
        RECT 394.185 50.825 394.565 51.205 ;
        RECT 404.470 50.825 404.850 51.205 ;
        RECT 414.760 50.825 415.140 51.205 ;
        RECT 425.045 50.825 425.425 51.205 ;
        RECT 426.465 50.825 426.845 51.205 ;
        RECT 436.755 50.825 437.135 51.205 ;
        RECT 447.040 50.825 447.420 51.205 ;
        RECT 457.330 50.825 457.710 51.205 ;
        RECT 467.615 50.825 467.995 51.205 ;
        RECT 469.035 50.825 469.415 51.205 ;
        RECT 479.325 50.825 479.705 51.205 ;
        RECT 489.610 50.825 489.990 51.205 ;
        RECT 499.900 50.825 500.280 51.205 ;
        RECT 510.185 50.825 510.565 51.205 ;
        RECT 511.605 50.825 511.985 51.205 ;
        RECT 521.895 50.825 522.275 51.205 ;
        RECT 532.180 50.825 532.560 51.205 ;
        RECT 542.470 50.825 542.850 51.205 ;
        RECT 552.755 50.825 553.135 51.205 ;
        RECT 554.175 50.825 554.555 51.205 ;
        RECT 564.465 50.825 564.845 51.205 ;
        RECT 574.750 50.825 575.130 51.205 ;
        RECT 585.040 50.825 585.420 51.205 ;
        RECT 595.325 50.825 595.705 51.205 ;
        RECT 596.745 50.825 597.125 51.205 ;
        RECT 607.035 50.825 607.415 51.205 ;
        RECT 617.320 50.825 617.700 51.205 ;
        RECT 627.610 50.825 627.990 51.205 ;
        RECT 637.895 50.825 638.275 51.205 ;
        RECT 639.315 50.825 639.695 51.205 ;
        RECT 649.605 50.825 649.985 51.205 ;
        RECT 659.890 50.825 660.270 51.205 ;
        RECT 670.180 50.825 670.560 51.205 ;
        RECT 680.465 50.825 680.845 51.205 ;
        RECT 682.310 51.155 682.690 51.535 ;
        RECT 684.095 51.155 684.475 51.535 ;
        RECT 686.950 51.155 687.330 51.535 ;
        RECT 688.735 51.155 689.115 51.535 ;
        RECT 691.590 51.155 691.970 51.535 ;
        RECT 693.375 51.155 693.755 51.535 ;
        RECT 696.230 51.155 696.610 51.535 ;
        RECT 698.015 51.155 698.395 51.535 ;
        RECT 700.870 51.155 701.250 51.535 ;
        RECT 702.655 51.155 703.035 51.535 ;
        RECT 705.510 51.155 705.890 51.535 ;
        RECT 707.295 51.155 707.675 51.535 ;
        RECT 710.150 51.155 710.530 51.535 ;
        RECT 711.935 51.155 712.315 51.535 ;
        RECT 714.790 51.155 715.170 51.535 ;
        RECT 716.575 51.155 716.955 51.535 ;
        RECT 0.765 50.165 1.145 50.545 ;
        RECT 11.055 50.165 11.435 50.545 ;
        RECT 21.340 50.165 21.720 50.545 ;
        RECT 31.630 50.165 32.010 50.545 ;
        RECT 41.915 50.165 42.295 50.545 ;
        RECT 43.335 50.165 43.715 50.545 ;
        RECT 53.625 50.165 54.005 50.545 ;
        RECT 63.910 50.165 64.290 50.545 ;
        RECT 74.200 50.165 74.580 50.545 ;
        RECT 84.485 50.165 84.865 50.545 ;
        RECT 85.905 50.165 86.285 50.545 ;
        RECT 96.195 50.165 96.575 50.545 ;
        RECT 106.480 50.165 106.860 50.545 ;
        RECT 116.770 50.165 117.150 50.545 ;
        RECT 127.055 50.165 127.435 50.545 ;
        RECT 128.475 50.165 128.855 50.545 ;
        RECT 138.765 50.165 139.145 50.545 ;
        RECT 149.050 50.165 149.430 50.545 ;
        RECT 159.340 50.165 159.720 50.545 ;
        RECT 169.625 50.165 170.005 50.545 ;
        RECT 171.045 50.165 171.425 50.545 ;
        RECT 181.335 50.165 181.715 50.545 ;
        RECT 191.620 50.165 192.000 50.545 ;
        RECT 201.910 50.165 202.290 50.545 ;
        RECT 212.195 50.165 212.575 50.545 ;
        RECT 213.615 50.165 213.995 50.545 ;
        RECT 223.905 50.165 224.285 50.545 ;
        RECT 234.190 50.165 234.570 50.545 ;
        RECT 244.480 50.165 244.860 50.545 ;
        RECT 254.765 50.165 255.145 50.545 ;
        RECT 256.185 50.165 256.565 50.545 ;
        RECT 266.475 50.165 266.855 50.545 ;
        RECT 276.760 50.165 277.140 50.545 ;
        RECT 287.050 50.165 287.430 50.545 ;
        RECT 297.335 50.165 297.715 50.545 ;
        RECT 298.755 50.165 299.135 50.545 ;
        RECT 309.045 50.165 309.425 50.545 ;
        RECT 319.330 50.165 319.710 50.545 ;
        RECT 329.620 50.165 330.000 50.545 ;
        RECT 339.905 50.165 340.285 50.545 ;
        RECT 341.325 50.165 341.705 50.545 ;
        RECT 351.615 50.165 351.995 50.545 ;
        RECT 361.900 50.165 362.280 50.545 ;
        RECT 372.190 50.165 372.570 50.545 ;
        RECT 382.475 50.165 382.855 50.545 ;
        RECT 383.895 50.165 384.275 50.545 ;
        RECT 394.185 50.165 394.565 50.545 ;
        RECT 404.470 50.165 404.850 50.545 ;
        RECT 414.760 50.165 415.140 50.545 ;
        RECT 425.045 50.165 425.425 50.545 ;
        RECT 426.465 50.165 426.845 50.545 ;
        RECT 436.755 50.165 437.135 50.545 ;
        RECT 447.040 50.165 447.420 50.545 ;
        RECT 457.330 50.165 457.710 50.545 ;
        RECT 467.615 50.165 467.995 50.545 ;
        RECT 469.035 50.165 469.415 50.545 ;
        RECT 479.325 50.165 479.705 50.545 ;
        RECT 489.610 50.165 489.990 50.545 ;
        RECT 499.900 50.165 500.280 50.545 ;
        RECT 510.185 50.165 510.565 50.545 ;
        RECT 511.605 50.165 511.985 50.545 ;
        RECT 521.895 50.165 522.275 50.545 ;
        RECT 532.180 50.165 532.560 50.545 ;
        RECT 542.470 50.165 542.850 50.545 ;
        RECT 552.755 50.165 553.135 50.545 ;
        RECT 554.175 50.165 554.555 50.545 ;
        RECT 564.465 50.165 564.845 50.545 ;
        RECT 574.750 50.165 575.130 50.545 ;
        RECT 585.040 50.165 585.420 50.545 ;
        RECT 595.325 50.165 595.705 50.545 ;
        RECT 596.745 50.165 597.125 50.545 ;
        RECT 607.035 50.165 607.415 50.545 ;
        RECT 617.320 50.165 617.700 50.545 ;
        RECT 627.610 50.165 627.990 50.545 ;
        RECT 637.895 50.165 638.275 50.545 ;
        RECT 639.315 50.165 639.695 50.545 ;
        RECT 649.605 50.165 649.985 50.545 ;
        RECT 659.890 50.165 660.270 50.545 ;
        RECT 670.180 50.165 670.560 50.545 ;
        RECT 680.465 50.165 680.845 50.545 ;
        RECT 682.310 50.495 682.690 50.875 ;
        RECT 684.095 50.495 684.475 50.875 ;
        RECT 686.950 50.495 687.330 50.875 ;
        RECT 688.735 50.495 689.115 50.875 ;
        RECT 691.590 50.495 691.970 50.875 ;
        RECT 693.375 50.495 693.755 50.875 ;
        RECT 696.230 50.495 696.610 50.875 ;
        RECT 698.015 50.495 698.395 50.875 ;
        RECT 700.870 50.495 701.250 50.875 ;
        RECT 702.655 50.495 703.035 50.875 ;
        RECT 705.510 50.495 705.890 50.875 ;
        RECT 707.295 50.495 707.675 50.875 ;
        RECT 710.150 50.495 710.530 50.875 ;
        RECT 711.935 50.495 712.315 50.875 ;
        RECT 714.790 50.495 715.170 50.875 ;
        RECT 716.575 50.495 716.955 50.875 ;
        RECT 0.500 46.485 717.540 48.185 ;
        RECT 0.500 43.785 717.540 45.485 ;
        RECT 0.500 41.085 717.540 42.785 ;
        RECT 0.500 38.385 717.540 40.085 ;
        RECT 0.500 28.985 717.540 30.685 ;
        RECT 0.500 26.285 717.540 27.985 ;
        RECT 0.500 23.585 717.540 25.285 ;
        RECT 0.500 20.885 717.540 22.585 ;
        RECT 682.310 18.115 682.690 18.495 ;
        RECT 684.095 18.115 684.475 18.495 ;
        RECT 686.950 18.115 687.330 18.495 ;
        RECT 688.735 18.115 689.115 18.495 ;
        RECT 691.590 18.115 691.970 18.495 ;
        RECT 693.375 18.115 693.755 18.495 ;
        RECT 696.230 18.115 696.610 18.495 ;
        RECT 698.015 18.115 698.395 18.495 ;
        RECT 700.870 18.115 701.250 18.495 ;
        RECT 702.655 18.115 703.035 18.495 ;
        RECT 705.510 18.115 705.890 18.495 ;
        RECT 707.295 18.115 707.675 18.495 ;
        RECT 710.150 18.115 710.530 18.495 ;
        RECT 711.935 18.115 712.315 18.495 ;
        RECT 714.790 18.115 715.170 18.495 ;
        RECT 716.575 18.115 716.955 18.495 ;
        RECT 682.310 17.455 682.690 17.835 ;
        RECT 684.095 17.455 684.475 17.835 ;
        RECT 686.950 17.455 687.330 17.835 ;
        RECT 688.735 17.455 689.115 17.835 ;
        RECT 691.590 17.455 691.970 17.835 ;
        RECT 693.375 17.455 693.755 17.835 ;
        RECT 696.230 17.455 696.610 17.835 ;
        RECT 698.015 17.455 698.395 17.835 ;
        RECT 700.870 17.455 701.250 17.835 ;
        RECT 702.655 17.455 703.035 17.835 ;
        RECT 705.510 17.455 705.890 17.835 ;
        RECT 707.295 17.455 707.675 17.835 ;
        RECT 710.150 17.455 710.530 17.835 ;
        RECT 711.935 17.455 712.315 17.835 ;
        RECT 714.790 17.455 715.170 17.835 ;
        RECT 716.575 17.455 716.955 17.835 ;
        RECT 682.310 16.795 682.690 17.175 ;
        RECT 684.095 16.795 684.475 17.175 ;
        RECT 686.950 16.795 687.330 17.175 ;
        RECT 688.735 16.795 689.115 17.175 ;
        RECT 691.590 16.795 691.970 17.175 ;
        RECT 693.375 16.795 693.755 17.175 ;
        RECT 696.230 16.795 696.610 17.175 ;
        RECT 698.015 16.795 698.395 17.175 ;
        RECT 700.870 16.795 701.250 17.175 ;
        RECT 702.655 16.795 703.035 17.175 ;
        RECT 705.510 16.795 705.890 17.175 ;
        RECT 707.295 16.795 707.675 17.175 ;
        RECT 710.150 16.795 710.530 17.175 ;
        RECT 711.935 16.795 712.315 17.175 ;
        RECT 714.790 16.795 715.170 17.175 ;
        RECT 716.575 16.795 716.955 17.175 ;
        RECT 682.310 16.135 682.690 16.515 ;
        RECT 684.095 16.135 684.475 16.515 ;
        RECT 686.950 16.135 687.330 16.515 ;
        RECT 688.735 16.135 689.115 16.515 ;
        RECT 691.590 16.135 691.970 16.515 ;
        RECT 693.375 16.135 693.755 16.515 ;
        RECT 696.230 16.135 696.610 16.515 ;
        RECT 698.015 16.135 698.395 16.515 ;
        RECT 700.870 16.135 701.250 16.515 ;
        RECT 702.655 16.135 703.035 16.515 ;
        RECT 705.510 16.135 705.890 16.515 ;
        RECT 707.295 16.135 707.675 16.515 ;
        RECT 710.150 16.135 710.530 16.515 ;
        RECT 711.935 16.135 712.315 16.515 ;
        RECT 714.790 16.135 715.170 16.515 ;
        RECT 716.575 16.135 716.955 16.515 ;
        RECT 682.310 15.475 682.690 15.855 ;
        RECT 684.095 15.475 684.475 15.855 ;
        RECT 686.950 15.475 687.330 15.855 ;
        RECT 688.735 15.475 689.115 15.855 ;
        RECT 691.590 15.475 691.970 15.855 ;
        RECT 693.375 15.475 693.755 15.855 ;
        RECT 696.230 15.475 696.610 15.855 ;
        RECT 698.015 15.475 698.395 15.855 ;
        RECT 700.870 15.475 701.250 15.855 ;
        RECT 702.655 15.475 703.035 15.855 ;
        RECT 705.510 15.475 705.890 15.855 ;
        RECT 707.295 15.475 707.675 15.855 ;
        RECT 710.150 15.475 710.530 15.855 ;
        RECT 711.935 15.475 712.315 15.855 ;
        RECT 714.790 15.475 715.170 15.855 ;
        RECT 716.575 15.475 716.955 15.855 ;
        RECT 682.310 14.815 682.690 15.195 ;
        RECT 684.095 14.815 684.475 15.195 ;
        RECT 686.950 14.815 687.330 15.195 ;
        RECT 688.735 14.815 689.115 15.195 ;
        RECT 691.590 14.815 691.970 15.195 ;
        RECT 693.375 14.815 693.755 15.195 ;
        RECT 696.230 14.815 696.610 15.195 ;
        RECT 698.015 14.815 698.395 15.195 ;
        RECT 700.870 14.815 701.250 15.195 ;
        RECT 702.655 14.815 703.035 15.195 ;
        RECT 705.510 14.815 705.890 15.195 ;
        RECT 707.295 14.815 707.675 15.195 ;
        RECT 710.150 14.815 710.530 15.195 ;
        RECT 711.935 14.815 712.315 15.195 ;
        RECT 714.790 14.815 715.170 15.195 ;
        RECT 716.575 14.815 716.955 15.195 ;
        RECT 682.310 14.155 682.690 14.535 ;
        RECT 684.095 14.155 684.475 14.535 ;
        RECT 686.950 14.155 687.330 14.535 ;
        RECT 688.735 14.155 689.115 14.535 ;
        RECT 691.590 14.155 691.970 14.535 ;
        RECT 693.375 14.155 693.755 14.535 ;
        RECT 696.230 14.155 696.610 14.535 ;
        RECT 698.015 14.155 698.395 14.535 ;
        RECT 700.870 14.155 701.250 14.535 ;
        RECT 702.655 14.155 703.035 14.535 ;
        RECT 705.510 14.155 705.890 14.535 ;
        RECT 707.295 14.155 707.675 14.535 ;
        RECT 710.150 14.155 710.530 14.535 ;
        RECT 711.935 14.155 712.315 14.535 ;
        RECT 714.790 14.155 715.170 14.535 ;
        RECT 716.575 14.155 716.955 14.535 ;
        RECT 682.310 13.495 682.690 13.875 ;
        RECT 684.095 13.495 684.475 13.875 ;
        RECT 686.950 13.495 687.330 13.875 ;
        RECT 688.735 13.495 689.115 13.875 ;
        RECT 691.590 13.495 691.970 13.875 ;
        RECT 693.375 13.495 693.755 13.875 ;
        RECT 696.230 13.495 696.610 13.875 ;
        RECT 698.015 13.495 698.395 13.875 ;
        RECT 700.870 13.495 701.250 13.875 ;
        RECT 702.655 13.495 703.035 13.875 ;
        RECT 705.510 13.495 705.890 13.875 ;
        RECT 707.295 13.495 707.675 13.875 ;
        RECT 710.150 13.495 710.530 13.875 ;
        RECT 711.935 13.495 712.315 13.875 ;
        RECT 714.790 13.495 715.170 13.875 ;
        RECT 716.575 13.495 716.955 13.875 ;
        RECT 682.310 12.835 682.690 13.215 ;
        RECT 684.095 12.835 684.475 13.215 ;
        RECT 686.950 12.835 687.330 13.215 ;
        RECT 688.735 12.835 689.115 13.215 ;
        RECT 691.590 12.835 691.970 13.215 ;
        RECT 693.375 12.835 693.755 13.215 ;
        RECT 696.230 12.835 696.610 13.215 ;
        RECT 698.015 12.835 698.395 13.215 ;
        RECT 700.870 12.835 701.250 13.215 ;
        RECT 702.655 12.835 703.035 13.215 ;
        RECT 705.510 12.835 705.890 13.215 ;
        RECT 707.295 12.835 707.675 13.215 ;
        RECT 710.150 12.835 710.530 13.215 ;
        RECT 711.935 12.835 712.315 13.215 ;
        RECT 714.790 12.835 715.170 13.215 ;
        RECT 716.575 12.835 716.955 13.215 ;
        RECT 682.310 12.175 682.690 12.555 ;
        RECT 684.095 12.175 684.475 12.555 ;
        RECT 686.950 12.175 687.330 12.555 ;
        RECT 688.735 12.175 689.115 12.555 ;
        RECT 691.590 12.175 691.970 12.555 ;
        RECT 693.375 12.175 693.755 12.555 ;
        RECT 696.230 12.175 696.610 12.555 ;
        RECT 698.015 12.175 698.395 12.555 ;
        RECT 700.870 12.175 701.250 12.555 ;
        RECT 702.655 12.175 703.035 12.555 ;
        RECT 705.510 12.175 705.890 12.555 ;
        RECT 707.295 12.175 707.675 12.555 ;
        RECT 710.150 12.175 710.530 12.555 ;
        RECT 711.935 12.175 712.315 12.555 ;
        RECT 714.790 12.175 715.170 12.555 ;
        RECT 716.575 12.175 716.955 12.555 ;
        RECT 682.310 11.515 682.690 11.895 ;
        RECT 684.095 11.515 684.475 11.895 ;
        RECT 686.950 11.515 687.330 11.895 ;
        RECT 688.735 11.515 689.115 11.895 ;
        RECT 691.590 11.515 691.970 11.895 ;
        RECT 693.375 11.515 693.755 11.895 ;
        RECT 696.230 11.515 696.610 11.895 ;
        RECT 698.015 11.515 698.395 11.895 ;
        RECT 700.870 11.515 701.250 11.895 ;
        RECT 702.655 11.515 703.035 11.895 ;
        RECT 705.510 11.515 705.890 11.895 ;
        RECT 707.295 11.515 707.675 11.895 ;
        RECT 710.150 11.515 710.530 11.895 ;
        RECT 711.935 11.515 712.315 11.895 ;
        RECT 714.790 11.515 715.170 11.895 ;
        RECT 716.575 11.515 716.955 11.895 ;
        RECT 682.310 10.855 682.690 11.235 ;
        RECT 684.095 10.855 684.475 11.235 ;
        RECT 686.950 10.855 687.330 11.235 ;
        RECT 688.735 10.855 689.115 11.235 ;
        RECT 691.590 10.855 691.970 11.235 ;
        RECT 693.375 10.855 693.755 11.235 ;
        RECT 696.230 10.855 696.610 11.235 ;
        RECT 698.015 10.855 698.395 11.235 ;
        RECT 700.870 10.855 701.250 11.235 ;
        RECT 702.655 10.855 703.035 11.235 ;
        RECT 705.510 10.855 705.890 11.235 ;
        RECT 707.295 10.855 707.675 11.235 ;
        RECT 710.150 10.855 710.530 11.235 ;
        RECT 711.935 10.855 712.315 11.235 ;
        RECT 714.790 10.855 715.170 11.235 ;
        RECT 716.575 10.855 716.955 11.235 ;
        RECT 682.310 10.195 682.690 10.575 ;
        RECT 684.095 10.195 684.475 10.575 ;
        RECT 686.950 10.195 687.330 10.575 ;
        RECT 688.735 10.195 689.115 10.575 ;
        RECT 691.590 10.195 691.970 10.575 ;
        RECT 693.375 10.195 693.755 10.575 ;
        RECT 696.230 10.195 696.610 10.575 ;
        RECT 698.015 10.195 698.395 10.575 ;
        RECT 700.870 10.195 701.250 10.575 ;
        RECT 702.655 10.195 703.035 10.575 ;
        RECT 705.510 10.195 705.890 10.575 ;
        RECT 707.295 10.195 707.675 10.575 ;
        RECT 710.150 10.195 710.530 10.575 ;
        RECT 711.935 10.195 712.315 10.575 ;
        RECT 714.790 10.195 715.170 10.575 ;
        RECT 716.575 10.195 716.955 10.575 ;
        RECT 682.310 9.535 682.690 9.915 ;
        RECT 684.095 9.535 684.475 9.915 ;
        RECT 686.950 9.535 687.330 9.915 ;
        RECT 688.735 9.535 689.115 9.915 ;
        RECT 691.590 9.535 691.970 9.915 ;
        RECT 693.375 9.535 693.755 9.915 ;
        RECT 696.230 9.535 696.610 9.915 ;
        RECT 698.015 9.535 698.395 9.915 ;
        RECT 700.870 9.535 701.250 9.915 ;
        RECT 702.655 9.535 703.035 9.915 ;
        RECT 705.510 9.535 705.890 9.915 ;
        RECT 707.295 9.535 707.675 9.915 ;
        RECT 710.150 9.535 710.530 9.915 ;
        RECT 711.935 9.535 712.315 9.915 ;
        RECT 714.790 9.535 715.170 9.915 ;
        RECT 716.575 9.535 716.955 9.915 ;
        RECT 682.310 8.875 682.690 9.255 ;
        RECT 684.095 8.875 684.475 9.255 ;
        RECT 686.950 8.875 687.330 9.255 ;
        RECT 688.735 8.875 689.115 9.255 ;
        RECT 691.590 8.875 691.970 9.255 ;
        RECT 693.375 8.875 693.755 9.255 ;
        RECT 696.230 8.875 696.610 9.255 ;
        RECT 698.015 8.875 698.395 9.255 ;
        RECT 700.870 8.875 701.250 9.255 ;
        RECT 702.655 8.875 703.035 9.255 ;
        RECT 705.510 8.875 705.890 9.255 ;
        RECT 707.295 8.875 707.675 9.255 ;
        RECT 710.150 8.875 710.530 9.255 ;
        RECT 711.935 8.875 712.315 9.255 ;
        RECT 714.790 8.875 715.170 9.255 ;
        RECT 716.575 8.875 716.955 9.255 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 38.750 8.090 39.130 8.470 ;
        RECT 53.580 8.090 53.960 8.470 ;
        RECT 72.890 8.090 73.270 8.470 ;
        RECT 87.720 8.090 88.100 8.470 ;
        RECT 107.030 8.090 107.410 8.470 ;
        RECT 121.860 8.090 122.240 8.470 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 38.750 7.430 39.130 7.810 ;
        RECT 53.580 7.430 53.960 7.810 ;
        RECT 72.890 7.430 73.270 7.810 ;
        RECT 87.720 7.430 88.100 7.810 ;
        RECT 107.030 7.430 107.410 7.810 ;
        RECT 121.860 7.430 122.240 7.810 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 38.750 6.770 39.130 7.150 ;
        RECT 53.580 6.770 53.960 7.150 ;
        RECT 72.890 6.770 73.270 7.150 ;
        RECT 87.720 6.770 88.100 7.150 ;
        RECT 107.030 6.770 107.410 7.150 ;
        RECT 121.860 6.770 122.240 7.150 ;
        RECT 0.850 4.690 1.230 5.070 ;
        RECT 1.990 4.690 2.370 5.070 ;
        RECT 8.030 4.720 8.410 5.100 ;
        RECT 8.690 4.720 9.070 5.100 ;
        RECT 9.350 4.720 9.730 5.100 ;
        RECT 14.560 4.690 14.940 5.070 ;
        RECT 15.220 4.690 15.600 5.070 ;
        RECT 15.880 4.690 16.260 5.070 ;
        RECT 17.920 4.690 18.300 5.070 ;
        RECT 18.580 4.690 18.960 5.070 ;
        RECT 19.240 4.690 19.620 5.070 ;
        RECT 26.220 4.720 26.600 5.100 ;
        RECT 26.880 4.720 27.260 5.100 ;
        RECT 27.540 4.720 27.920 5.100 ;
        RECT 32.750 4.690 33.130 5.070 ;
        RECT 33.410 4.690 33.790 5.070 ;
        RECT 34.070 4.690 34.450 5.070 ;
        RECT 36.130 4.690 36.510 5.070 ;
        RECT 42.170 4.720 42.550 5.100 ;
        RECT 42.830 4.720 43.210 5.100 ;
        RECT 43.490 4.720 43.870 5.100 ;
        RECT 48.700 4.690 49.080 5.070 ;
        RECT 49.360 4.690 49.740 5.070 ;
        RECT 50.020 4.690 50.400 5.070 ;
        RECT 57.000 4.720 57.380 5.100 ;
        RECT 57.660 4.720 58.040 5.100 ;
        RECT 58.320 4.720 58.700 5.100 ;
        RECT 63.530 4.690 63.910 5.070 ;
        RECT 64.190 4.690 64.570 5.070 ;
        RECT 64.850 4.690 65.230 5.070 ;
        RECT 66.890 4.690 67.270 5.070 ;
        RECT 67.550 4.690 67.930 5.070 ;
        RECT 68.210 4.690 68.590 5.070 ;
        RECT 70.270 4.690 70.650 5.070 ;
        RECT 76.310 4.720 76.690 5.100 ;
        RECT 76.970 4.720 77.350 5.100 ;
        RECT 77.630 4.720 78.010 5.100 ;
        RECT 82.840 4.690 83.220 5.070 ;
        RECT 83.500 4.690 83.880 5.070 ;
        RECT 84.160 4.690 84.540 5.070 ;
        RECT 91.140 4.720 91.520 5.100 ;
        RECT 91.800 4.720 92.180 5.100 ;
        RECT 92.460 4.720 92.840 5.100 ;
        RECT 97.670 4.690 98.050 5.070 ;
        RECT 98.330 4.690 98.710 5.070 ;
        RECT 98.990 4.690 99.370 5.070 ;
        RECT 101.030 4.690 101.410 5.070 ;
        RECT 101.690 4.690 102.070 5.070 ;
        RECT 102.350 4.690 102.730 5.070 ;
        RECT 104.410 4.690 104.790 5.070 ;
        RECT 110.450 4.720 110.830 5.100 ;
        RECT 111.110 4.720 111.490 5.100 ;
        RECT 111.770 4.720 112.150 5.100 ;
        RECT 116.980 4.690 117.360 5.070 ;
        RECT 117.640 4.690 118.020 5.070 ;
        RECT 118.300 4.690 118.680 5.070 ;
        RECT 125.280 4.720 125.660 5.100 ;
        RECT 125.940 4.720 126.320 5.100 ;
        RECT 126.600 4.720 126.980 5.100 ;
        RECT 131.810 4.690 132.190 5.070 ;
        RECT 132.470 4.690 132.850 5.070 ;
        RECT 133.130 4.690 133.510 5.070 ;
        RECT 135.190 4.690 135.570 5.070 ;
        RECT 136.190 4.690 136.570 5.070 ;
        RECT 136.850 4.690 137.230 5.070 ;
        RECT 137.510 4.690 137.890 5.070 ;
        RECT 138.430 4.690 138.810 5.070 ;
        RECT 139.090 4.690 139.470 5.070 ;
        RECT 139.750 4.690 140.130 5.070 ;
        RECT 140.770 4.690 141.150 5.070 ;
        RECT 141.430 4.690 141.810 5.070 ;
        RECT 142.090 4.690 142.470 5.070 ;
        RECT 144.030 4.690 144.410 5.070 ;
        RECT 144.690 4.690 145.070 5.070 ;
        RECT 145.350 4.690 145.730 5.070 ;
        RECT 146.270 4.690 146.650 5.070 ;
        RECT 146.930 4.690 147.310 5.070 ;
        RECT 147.590 4.690 147.970 5.070 ;
        RECT 148.510 4.690 148.890 5.070 ;
        RECT 149.170 4.690 149.550 5.070 ;
        RECT 149.830 4.690 150.210 5.070 ;
        RECT 150.750 4.690 151.130 5.070 ;
        RECT 151.410 4.690 151.790 5.070 ;
        RECT 152.070 4.690 152.450 5.070 ;
        RECT 152.990 4.690 153.370 5.070 ;
        RECT 153.650 4.690 154.030 5.070 ;
        RECT 154.310 4.690 154.690 5.070 ;
        RECT 155.350 4.690 155.730 5.070 ;
        RECT 156.350 4.690 156.730 5.070 ;
        RECT 157.010 4.690 157.390 5.070 ;
        RECT 157.670 4.690 158.050 5.070 ;
        RECT 158.590 4.690 158.970 5.070 ;
        RECT 159.250 4.690 159.630 5.070 ;
        RECT 159.910 4.690 160.290 5.070 ;
        RECT 160.830 4.690 161.210 5.070 ;
        RECT 161.490 4.690 161.870 5.070 ;
        RECT 162.150 4.690 162.530 5.070 ;
        RECT 163.070 4.690 163.450 5.070 ;
        RECT 163.730 4.690 164.110 5.070 ;
        RECT 164.390 4.690 164.770 5.070 ;
        RECT 165.310 4.690 165.690 5.070 ;
        RECT 165.970 4.690 166.350 5.070 ;
        RECT 166.630 4.690 167.010 5.070 ;
        RECT 167.550 4.690 167.930 5.070 ;
        RECT 168.210 4.690 168.590 5.070 ;
        RECT 168.870 4.690 169.250 5.070 ;
        RECT 169.790 4.690 170.170 5.070 ;
        RECT 170.450 4.690 170.830 5.070 ;
        RECT 171.110 4.690 171.490 5.070 ;
        RECT 172.030 4.690 172.410 5.070 ;
        RECT 172.690 4.690 173.070 5.070 ;
        RECT 173.350 4.690 173.730 5.070 ;
        RECT 174.270 4.690 174.650 5.070 ;
        RECT 174.930 4.690 175.310 5.070 ;
        RECT 175.590 4.690 175.970 5.070 ;
        RECT 176.630 4.690 177.010 5.070 ;
        RECT 177.630 4.690 178.010 5.070 ;
        RECT 178.290 4.690 178.670 5.070 ;
        RECT 178.950 4.690 179.330 5.070 ;
        RECT 179.870 4.690 180.250 5.070 ;
        RECT 180.530 4.690 180.910 5.070 ;
        RECT 181.190 4.690 181.570 5.070 ;
        RECT 182.210 4.690 182.590 5.070 ;
        RECT 182.870 4.690 183.250 5.070 ;
        RECT 183.530 4.690 183.910 5.070 ;
        RECT 185.470 4.690 185.850 5.070 ;
        RECT 186.130 4.690 186.510 5.070 ;
        RECT 186.790 4.690 187.170 5.070 ;
        RECT 187.710 4.690 188.090 5.070 ;
        RECT 188.370 4.690 188.750 5.070 ;
        RECT 189.030 4.690 189.410 5.070 ;
        RECT 189.950 4.690 190.330 5.070 ;
        RECT 190.610 4.690 190.990 5.070 ;
        RECT 191.270 4.690 191.650 5.070 ;
        RECT 192.190 4.690 192.570 5.070 ;
        RECT 192.850 4.690 193.230 5.070 ;
        RECT 193.510 4.690 193.890 5.070 ;
        RECT 194.430 4.690 194.810 5.070 ;
        RECT 195.090 4.690 195.470 5.070 ;
        RECT 195.750 4.690 196.130 5.070 ;
        RECT 196.790 4.690 197.170 5.070 ;
        RECT 197.790 4.690 198.170 5.070 ;
        RECT 198.450 4.690 198.830 5.070 ;
        RECT 199.110 4.690 199.490 5.070 ;
        RECT 200.030 4.690 200.410 5.070 ;
        RECT 200.690 4.690 201.070 5.070 ;
        RECT 201.350 4.690 201.730 5.070 ;
        RECT 202.270 4.690 202.650 5.070 ;
        RECT 202.930 4.690 203.310 5.070 ;
        RECT 203.590 4.690 203.970 5.070 ;
        RECT 204.510 4.690 204.890 5.070 ;
        RECT 205.170 4.690 205.550 5.070 ;
        RECT 205.830 4.690 206.210 5.070 ;
        RECT 206.750 4.690 207.130 5.070 ;
        RECT 207.410 4.690 207.790 5.070 ;
        RECT 208.070 4.690 208.450 5.070 ;
        RECT 208.990 4.690 209.370 5.070 ;
        RECT 209.650 4.690 210.030 5.070 ;
        RECT 210.310 4.690 210.690 5.070 ;
        RECT 211.230 4.690 211.610 5.070 ;
        RECT 211.890 4.690 212.270 5.070 ;
        RECT 212.550 4.690 212.930 5.070 ;
        RECT 213.470 4.690 213.850 5.070 ;
        RECT 214.130 4.690 214.510 5.070 ;
        RECT 214.790 4.690 215.170 5.070 ;
        RECT 215.710 4.690 216.090 5.070 ;
        RECT 216.370 4.690 216.750 5.070 ;
        RECT 217.030 4.690 217.410 5.070 ;
        RECT 218.070 4.690 218.450 5.070 ;
        RECT 219.070 4.690 219.450 5.070 ;
        RECT 219.730 4.690 220.110 5.070 ;
        RECT 220.390 4.690 220.770 5.070 ;
        RECT 221.310 4.690 221.690 5.070 ;
        RECT 221.970 4.690 222.350 5.070 ;
        RECT 222.630 4.690 223.010 5.070 ;
        RECT 223.550 4.690 223.930 5.070 ;
        RECT 224.210 4.690 224.590 5.070 ;
        RECT 224.870 4.690 225.250 5.070 ;
        RECT 225.890 4.690 226.270 5.070 ;
        RECT 226.550 4.690 226.930 5.070 ;
        RECT 227.210 4.690 227.590 5.070 ;
        RECT 229.150 4.690 229.530 5.070 ;
        RECT 229.810 4.690 230.190 5.070 ;
        RECT 230.470 4.690 230.850 5.070 ;
        RECT 231.390 4.690 231.770 5.070 ;
        RECT 232.050 4.690 232.430 5.070 ;
        RECT 232.710 4.690 233.090 5.070 ;
        RECT 233.630 4.690 234.010 5.070 ;
        RECT 234.290 4.690 234.670 5.070 ;
        RECT 234.950 4.690 235.330 5.070 ;
        RECT 235.870 4.690 236.250 5.070 ;
        RECT 236.530 4.690 236.910 5.070 ;
        RECT 237.190 4.690 237.570 5.070 ;
        RECT 238.230 4.690 238.610 5.070 ;
        RECT 239.230 4.690 239.610 5.070 ;
        RECT 239.890 4.690 240.270 5.070 ;
        RECT 240.550 4.690 240.930 5.070 ;
        RECT 241.470 4.690 241.850 5.070 ;
        RECT 242.130 4.690 242.510 5.070 ;
        RECT 242.790 4.690 243.170 5.070 ;
        RECT 243.710 4.690 244.090 5.070 ;
        RECT 244.370 4.690 244.750 5.070 ;
        RECT 245.030 4.690 245.410 5.070 ;
        RECT 245.950 4.690 246.330 5.070 ;
        RECT 246.610 4.690 246.990 5.070 ;
        RECT 247.270 4.690 247.650 5.070 ;
        RECT 248.190 4.690 248.570 5.070 ;
        RECT 248.850 4.690 249.230 5.070 ;
        RECT 249.510 4.690 249.890 5.070 ;
        RECT 250.430 4.690 250.810 5.070 ;
        RECT 251.090 4.690 251.470 5.070 ;
        RECT 251.750 4.690 252.130 5.070 ;
        RECT 252.670 4.690 253.050 5.070 ;
        RECT 253.330 4.690 253.710 5.070 ;
        RECT 253.990 4.690 254.370 5.070 ;
        RECT 254.910 4.690 255.290 5.070 ;
        RECT 255.570 4.690 255.950 5.070 ;
        RECT 256.230 4.690 256.610 5.070 ;
        RECT 257.150 4.690 257.530 5.070 ;
        RECT 257.810 4.690 258.190 5.070 ;
        RECT 258.470 4.690 258.850 5.070 ;
        RECT 259.510 4.690 259.890 5.070 ;
        RECT 260.510 4.690 260.890 5.070 ;
        RECT 261.170 4.690 261.550 5.070 ;
        RECT 261.830 4.690 262.210 5.070 ;
        RECT 262.750 4.690 263.130 5.070 ;
        RECT 263.410 4.690 263.790 5.070 ;
        RECT 264.070 4.690 264.450 5.070 ;
        RECT 264.990 4.690 265.370 5.070 ;
        RECT 265.650 4.690 266.030 5.070 ;
        RECT 266.310 4.690 266.690 5.070 ;
        RECT 267.330 4.690 267.710 5.070 ;
        RECT 267.990 4.690 268.370 5.070 ;
        RECT 268.650 4.690 269.030 5.070 ;
        RECT 270.590 4.690 270.970 5.070 ;
        RECT 271.250 4.690 271.630 5.070 ;
        RECT 271.910 4.690 272.290 5.070 ;
        RECT 272.830 4.690 273.210 5.070 ;
        RECT 273.490 4.690 273.870 5.070 ;
        RECT 274.150 4.690 274.530 5.070 ;
        RECT 275.070 4.690 275.450 5.070 ;
        RECT 275.730 4.690 276.110 5.070 ;
        RECT 276.390 4.690 276.770 5.070 ;
        RECT 277.310 4.690 277.690 5.070 ;
        RECT 277.970 4.690 278.350 5.070 ;
        RECT 278.630 4.690 279.010 5.070 ;
        RECT 279.670 4.690 280.050 5.070 ;
        RECT 280.670 4.690 281.050 5.070 ;
        RECT 281.330 4.690 281.710 5.070 ;
        RECT 281.990 4.690 282.370 5.070 ;
        RECT 282.910 4.690 283.290 5.070 ;
        RECT 283.570 4.690 283.950 5.070 ;
        RECT 284.230 4.690 284.610 5.070 ;
        RECT 285.150 4.690 285.530 5.070 ;
        RECT 285.810 4.690 286.190 5.070 ;
        RECT 286.470 4.690 286.850 5.070 ;
        RECT 287.390 4.690 287.770 5.070 ;
        RECT 288.050 4.690 288.430 5.070 ;
        RECT 288.710 4.690 289.090 5.070 ;
        RECT 289.630 4.690 290.010 5.070 ;
        RECT 290.290 4.690 290.670 5.070 ;
        RECT 290.950 4.690 291.330 5.070 ;
        RECT 291.870 4.690 292.250 5.070 ;
        RECT 292.530 4.690 292.910 5.070 ;
        RECT 293.190 4.690 293.570 5.070 ;
        RECT 294.110 4.690 294.490 5.070 ;
        RECT 294.770 4.690 295.150 5.070 ;
        RECT 295.430 4.690 295.810 5.070 ;
        RECT 296.350 4.690 296.730 5.070 ;
        RECT 297.010 4.690 297.390 5.070 ;
        RECT 297.670 4.690 298.050 5.070 ;
        RECT 298.590 4.690 298.970 5.070 ;
        RECT 299.250 4.690 299.630 5.070 ;
        RECT 299.910 4.690 300.290 5.070 ;
        RECT 300.950 4.690 301.330 5.070 ;
        RECT 301.950 4.690 302.330 5.070 ;
        RECT 302.610 4.690 302.990 5.070 ;
        RECT 303.270 4.690 303.650 5.070 ;
        RECT 304.190 4.690 304.570 5.070 ;
        RECT 304.850 4.690 305.230 5.070 ;
        RECT 305.510 4.690 305.890 5.070 ;
        RECT 306.430 4.690 306.810 5.070 ;
        RECT 307.090 4.690 307.470 5.070 ;
        RECT 307.750 4.690 308.130 5.070 ;
        RECT 308.670 4.690 309.050 5.070 ;
        RECT 309.330 4.690 309.710 5.070 ;
        RECT 309.990 4.690 310.370 5.070 ;
        RECT 311.010 4.690 311.390 5.070 ;
        RECT 311.670 4.690 312.050 5.070 ;
        RECT 312.330 4.690 312.710 5.070 ;
        RECT 314.270 4.690 314.650 5.070 ;
        RECT 314.930 4.690 315.310 5.070 ;
        RECT 315.590 4.690 315.970 5.070 ;
        RECT 316.510 4.690 316.890 5.070 ;
        RECT 317.170 4.690 317.550 5.070 ;
        RECT 317.830 4.690 318.210 5.070 ;
        RECT 318.750 4.690 319.130 5.070 ;
        RECT 319.410 4.690 319.790 5.070 ;
        RECT 320.070 4.690 320.450 5.070 ;
        RECT 321.110 4.690 321.490 5.070 ;
        RECT 322.110 4.690 322.490 5.070 ;
        RECT 322.770 4.690 323.150 5.070 ;
        RECT 323.430 4.690 323.810 5.070 ;
        RECT 324.350 4.690 324.730 5.070 ;
        RECT 325.010 4.690 325.390 5.070 ;
        RECT 325.670 4.690 326.050 5.070 ;
        RECT 326.590 4.690 326.970 5.070 ;
        RECT 327.250 4.690 327.630 5.070 ;
        RECT 327.910 4.690 328.290 5.070 ;
        RECT 328.830 4.690 329.210 5.070 ;
        RECT 329.490 4.690 329.870 5.070 ;
        RECT 330.150 4.690 330.530 5.070 ;
        RECT 331.070 4.690 331.450 5.070 ;
        RECT 331.730 4.690 332.110 5.070 ;
        RECT 332.390 4.690 332.770 5.070 ;
        RECT 333.310 4.690 333.690 5.070 ;
        RECT 333.970 4.690 334.350 5.070 ;
        RECT 334.630 4.690 335.010 5.070 ;
        RECT 335.550 4.690 335.930 5.070 ;
        RECT 336.210 4.690 336.590 5.070 ;
        RECT 336.870 4.690 337.250 5.070 ;
        RECT 337.790 4.690 338.170 5.070 ;
        RECT 338.450 4.690 338.830 5.070 ;
        RECT 339.110 4.690 339.490 5.070 ;
        RECT 340.030 4.690 340.410 5.070 ;
        RECT 340.690 4.690 341.070 5.070 ;
        RECT 341.350 4.690 341.730 5.070 ;
        RECT 342.390 4.690 342.770 5.070 ;
        RECT 343.390 4.690 343.770 5.070 ;
        RECT 344.050 4.690 344.430 5.070 ;
        RECT 344.710 4.690 345.090 5.070 ;
        RECT 345.630 4.690 346.010 5.070 ;
        RECT 346.290 4.690 346.670 5.070 ;
        RECT 346.950 4.690 347.330 5.070 ;
        RECT 347.870 4.690 348.250 5.070 ;
        RECT 348.530 4.690 348.910 5.070 ;
        RECT 349.190 4.690 349.570 5.070 ;
        RECT 350.110 4.690 350.490 5.070 ;
        RECT 350.770 4.690 351.150 5.070 ;
        RECT 351.430 4.690 351.810 5.070 ;
        RECT 352.450 4.690 352.830 5.070 ;
        RECT 353.110 4.690 353.490 5.070 ;
        RECT 353.770 4.690 354.150 5.070 ;
        RECT 355.710 4.690 356.090 5.070 ;
        RECT 356.370 4.690 356.750 5.070 ;
        RECT 357.030 4.690 357.410 5.070 ;
        RECT 357.950 4.690 358.330 5.070 ;
        RECT 358.610 4.690 358.990 5.070 ;
        RECT 359.270 4.690 359.650 5.070 ;
        RECT 360.190 4.690 360.570 5.070 ;
        RECT 360.850 4.690 361.230 5.070 ;
        RECT 361.510 4.690 361.890 5.070 ;
        RECT 362.550 4.690 362.930 5.070 ;
        RECT 363.550 4.690 363.930 5.070 ;
        RECT 364.210 4.690 364.590 5.070 ;
        RECT 364.870 4.690 365.250 5.070 ;
        RECT 365.790 4.690 366.170 5.070 ;
        RECT 366.450 4.690 366.830 5.070 ;
        RECT 367.110 4.690 367.490 5.070 ;
        RECT 368.030 4.690 368.410 5.070 ;
        RECT 368.690 4.690 369.070 5.070 ;
        RECT 369.350 4.690 369.730 5.070 ;
        RECT 370.270 4.690 370.650 5.070 ;
        RECT 370.930 4.690 371.310 5.070 ;
        RECT 371.590 4.690 371.970 5.070 ;
        RECT 372.510 4.690 372.890 5.070 ;
        RECT 373.170 4.690 373.550 5.070 ;
        RECT 373.830 4.690 374.210 5.070 ;
        RECT 374.750 4.690 375.130 5.070 ;
        RECT 375.410 4.690 375.790 5.070 ;
        RECT 376.070 4.690 376.450 5.070 ;
        RECT 376.990 4.690 377.370 5.070 ;
        RECT 377.650 4.690 378.030 5.070 ;
        RECT 378.310 4.690 378.690 5.070 ;
        RECT 379.230 4.690 379.610 5.070 ;
        RECT 379.890 4.690 380.270 5.070 ;
        RECT 380.550 4.690 380.930 5.070 ;
        RECT 381.470 4.690 381.850 5.070 ;
        RECT 382.130 4.690 382.510 5.070 ;
        RECT 382.790 4.690 383.170 5.070 ;
        RECT 383.830 4.690 384.210 5.070 ;
        RECT 384.830 4.690 385.210 5.070 ;
        RECT 385.490 4.690 385.870 5.070 ;
        RECT 386.150 4.690 386.530 5.070 ;
        RECT 387.070 4.690 387.450 5.070 ;
        RECT 387.730 4.690 388.110 5.070 ;
        RECT 388.390 4.690 388.770 5.070 ;
        RECT 389.310 4.690 389.690 5.070 ;
        RECT 389.970 4.690 390.350 5.070 ;
        RECT 390.630 4.690 391.010 5.070 ;
        RECT 391.550 4.690 391.930 5.070 ;
        RECT 392.210 4.690 392.590 5.070 ;
        RECT 392.870 4.690 393.250 5.070 ;
        RECT 393.790 4.690 394.170 5.070 ;
        RECT 394.450 4.690 394.830 5.070 ;
        RECT 395.110 4.690 395.490 5.070 ;
        RECT 396.130 4.690 396.510 5.070 ;
        RECT 396.790 4.690 397.170 5.070 ;
        RECT 397.450 4.690 397.830 5.070 ;
        RECT 399.390 4.690 399.770 5.070 ;
        RECT 400.050 4.690 400.430 5.070 ;
        RECT 400.710 4.690 401.090 5.070 ;
        RECT 401.630 4.690 402.010 5.070 ;
        RECT 402.290 4.690 402.670 5.070 ;
        RECT 402.950 4.690 403.330 5.070 ;
        RECT 403.990 4.690 404.370 5.070 ;
        RECT 404.990 4.690 405.370 5.070 ;
        RECT 405.650 4.690 406.030 5.070 ;
        RECT 406.310 4.690 406.690 5.070 ;
        RECT 407.230 4.690 407.610 5.070 ;
        RECT 407.890 4.690 408.270 5.070 ;
        RECT 408.550 4.690 408.930 5.070 ;
        RECT 409.470 4.690 409.850 5.070 ;
        RECT 410.130 4.690 410.510 5.070 ;
        RECT 410.790 4.690 411.170 5.070 ;
        RECT 411.710 4.690 412.090 5.070 ;
        RECT 412.370 4.690 412.750 5.070 ;
        RECT 413.030 4.690 413.410 5.070 ;
        RECT 413.950 4.690 414.330 5.070 ;
        RECT 414.610 4.690 414.990 5.070 ;
        RECT 415.270 4.690 415.650 5.070 ;
        RECT 416.190 4.690 416.570 5.070 ;
        RECT 416.850 4.690 417.230 5.070 ;
        RECT 417.510 4.690 417.890 5.070 ;
        RECT 418.430 4.690 418.810 5.070 ;
        RECT 419.090 4.690 419.470 5.070 ;
        RECT 419.750 4.690 420.130 5.070 ;
        RECT 420.670 4.690 421.050 5.070 ;
        RECT 421.330 4.690 421.710 5.070 ;
        RECT 421.990 4.690 422.370 5.070 ;
        RECT 422.910 4.690 423.290 5.070 ;
        RECT 423.570 4.690 423.950 5.070 ;
        RECT 424.230 4.690 424.610 5.070 ;
        RECT 425.270 4.690 425.650 5.070 ;
        RECT 426.270 4.690 426.650 5.070 ;
        RECT 426.930 4.690 427.310 5.070 ;
        RECT 427.590 4.690 427.970 5.070 ;
        RECT 428.510 4.690 428.890 5.070 ;
        RECT 429.170 4.690 429.550 5.070 ;
        RECT 429.830 4.690 430.210 5.070 ;
        RECT 430.750 4.690 431.130 5.070 ;
        RECT 431.410 4.690 431.790 5.070 ;
        RECT 432.070 4.690 432.450 5.070 ;
        RECT 432.990 4.690 433.370 5.070 ;
        RECT 433.650 4.690 434.030 5.070 ;
        RECT 434.310 4.690 434.690 5.070 ;
        RECT 435.230 4.690 435.610 5.070 ;
        RECT 435.890 4.690 436.270 5.070 ;
        RECT 436.550 4.690 436.930 5.070 ;
        RECT 437.570 4.690 437.950 5.070 ;
        RECT 438.230 4.690 438.610 5.070 ;
        RECT 438.890 4.690 439.270 5.070 ;
        RECT 440.830 4.690 441.210 5.070 ;
        RECT 441.490 4.690 441.870 5.070 ;
        RECT 442.150 4.690 442.530 5.070 ;
        RECT 443.070 4.690 443.450 5.070 ;
        RECT 443.730 4.690 444.110 5.070 ;
        RECT 444.390 4.690 444.770 5.070 ;
        RECT 445.430 4.690 445.810 5.070 ;
        RECT 446.430 4.690 446.810 5.070 ;
        RECT 447.090 4.690 447.470 5.070 ;
        RECT 447.750 4.690 448.130 5.070 ;
        RECT 448.670 4.690 449.050 5.070 ;
        RECT 449.330 4.690 449.710 5.070 ;
        RECT 449.990 4.690 450.370 5.070 ;
        RECT 450.910 4.690 451.290 5.070 ;
        RECT 451.570 4.690 451.950 5.070 ;
        RECT 452.230 4.690 452.610 5.070 ;
        RECT 453.150 4.690 453.530 5.070 ;
        RECT 453.810 4.690 454.190 5.070 ;
        RECT 454.470 4.690 454.850 5.070 ;
        RECT 455.390 4.690 455.770 5.070 ;
        RECT 456.050 4.690 456.430 5.070 ;
        RECT 456.710 4.690 457.090 5.070 ;
        RECT 457.630 4.690 458.010 5.070 ;
        RECT 458.290 4.690 458.670 5.070 ;
        RECT 458.950 4.690 459.330 5.070 ;
        RECT 459.870 4.690 460.250 5.070 ;
        RECT 460.530 4.690 460.910 5.070 ;
        RECT 461.190 4.690 461.570 5.070 ;
        RECT 462.110 4.690 462.490 5.070 ;
        RECT 462.770 4.690 463.150 5.070 ;
        RECT 463.430 4.690 463.810 5.070 ;
        RECT 464.350 4.690 464.730 5.070 ;
        RECT 465.010 4.690 465.390 5.070 ;
        RECT 465.670 4.690 466.050 5.070 ;
        RECT 466.710 4.690 467.090 5.070 ;
        RECT 467.710 4.690 468.090 5.070 ;
        RECT 468.370 4.690 468.750 5.070 ;
        RECT 469.030 4.690 469.410 5.070 ;
        RECT 469.950 4.690 470.330 5.070 ;
        RECT 470.610 4.690 470.990 5.070 ;
        RECT 471.270 4.690 471.650 5.070 ;
        RECT 472.190 4.690 472.570 5.070 ;
        RECT 472.850 4.690 473.230 5.070 ;
        RECT 473.510 4.690 473.890 5.070 ;
        RECT 474.430 4.690 474.810 5.070 ;
        RECT 475.090 4.690 475.470 5.070 ;
        RECT 475.750 4.690 476.130 5.070 ;
        RECT 476.670 4.690 477.050 5.070 ;
        RECT 477.330 4.690 477.710 5.070 ;
        RECT 477.990 4.690 478.370 5.070 ;
        RECT 478.910 4.690 479.290 5.070 ;
        RECT 479.570 4.690 479.950 5.070 ;
        RECT 480.230 4.690 480.610 5.070 ;
        RECT 481.250 4.690 481.630 5.070 ;
        RECT 481.910 4.690 482.290 5.070 ;
        RECT 482.570 4.690 482.950 5.070 ;
        RECT 484.510 4.690 484.890 5.070 ;
        RECT 485.170 4.690 485.550 5.070 ;
        RECT 485.830 4.690 486.210 5.070 ;
        RECT 486.870 4.690 487.250 5.070 ;
        RECT 487.870 4.690 488.250 5.070 ;
        RECT 488.530 4.690 488.910 5.070 ;
        RECT 489.190 4.690 489.570 5.070 ;
        RECT 490.110 4.690 490.490 5.070 ;
        RECT 490.770 4.690 491.150 5.070 ;
        RECT 491.430 4.690 491.810 5.070 ;
        RECT 492.350 4.690 492.730 5.070 ;
        RECT 493.010 4.690 493.390 5.070 ;
        RECT 493.670 4.690 494.050 5.070 ;
        RECT 494.590 4.690 494.970 5.070 ;
        RECT 495.250 4.690 495.630 5.070 ;
        RECT 495.910 4.690 496.290 5.070 ;
        RECT 496.830 4.690 497.210 5.070 ;
        RECT 497.490 4.690 497.870 5.070 ;
        RECT 498.150 4.690 498.530 5.070 ;
        RECT 499.070 4.690 499.450 5.070 ;
        RECT 499.730 4.690 500.110 5.070 ;
        RECT 500.390 4.690 500.770 5.070 ;
        RECT 501.310 4.690 501.690 5.070 ;
        RECT 501.970 4.690 502.350 5.070 ;
        RECT 502.630 4.690 503.010 5.070 ;
        RECT 503.550 4.690 503.930 5.070 ;
        RECT 504.210 4.690 504.590 5.070 ;
        RECT 504.870 4.690 505.250 5.070 ;
        RECT 505.790 4.690 506.170 5.070 ;
        RECT 506.450 4.690 506.830 5.070 ;
        RECT 507.110 4.690 507.490 5.070 ;
        RECT 508.150 4.690 508.530 5.070 ;
        RECT 509.150 4.690 509.530 5.070 ;
        RECT 509.810 4.690 510.190 5.070 ;
        RECT 510.470 4.690 510.850 5.070 ;
        RECT 511.390 4.690 511.770 5.070 ;
        RECT 512.050 4.690 512.430 5.070 ;
        RECT 512.710 4.690 513.090 5.070 ;
        RECT 513.630 4.690 514.010 5.070 ;
        RECT 514.290 4.690 514.670 5.070 ;
        RECT 514.950 4.690 515.330 5.070 ;
        RECT 515.870 4.690 516.250 5.070 ;
        RECT 516.530 4.690 516.910 5.070 ;
        RECT 517.190 4.690 517.570 5.070 ;
        RECT 518.110 4.690 518.490 5.070 ;
        RECT 518.770 4.690 519.150 5.070 ;
        RECT 519.430 4.690 519.810 5.070 ;
        RECT 520.350 4.690 520.730 5.070 ;
        RECT 521.010 4.690 521.390 5.070 ;
        RECT 521.670 4.690 522.050 5.070 ;
        RECT 522.690 4.690 523.070 5.070 ;
        RECT 523.350 4.690 523.730 5.070 ;
        RECT 524.010 4.690 524.390 5.070 ;
        RECT 525.950 4.690 526.330 5.070 ;
        RECT 526.610 4.690 526.990 5.070 ;
        RECT 527.270 4.690 527.650 5.070 ;
        RECT 528.310 4.690 528.690 5.070 ;
        RECT 529.310 4.690 529.690 5.070 ;
        RECT 529.970 4.690 530.350 5.070 ;
        RECT 530.630 4.690 531.010 5.070 ;
        RECT 531.550 4.690 531.930 5.070 ;
        RECT 532.210 4.690 532.590 5.070 ;
        RECT 532.870 4.690 533.250 5.070 ;
        RECT 533.790 4.690 534.170 5.070 ;
        RECT 534.450 4.690 534.830 5.070 ;
        RECT 535.110 4.690 535.490 5.070 ;
        RECT 536.030 4.690 536.410 5.070 ;
        RECT 536.690 4.690 537.070 5.070 ;
        RECT 537.350 4.690 537.730 5.070 ;
        RECT 538.270 4.690 538.650 5.070 ;
        RECT 538.930 4.690 539.310 5.070 ;
        RECT 539.590 4.690 539.970 5.070 ;
        RECT 540.510 4.690 540.890 5.070 ;
        RECT 541.170 4.690 541.550 5.070 ;
        RECT 541.830 4.690 542.210 5.070 ;
        RECT 542.750 4.690 543.130 5.070 ;
        RECT 543.410 4.690 543.790 5.070 ;
        RECT 544.070 4.690 544.450 5.070 ;
        RECT 544.990 4.690 545.370 5.070 ;
        RECT 545.650 4.690 546.030 5.070 ;
        RECT 546.310 4.690 546.690 5.070 ;
        RECT 547.230 4.690 547.610 5.070 ;
        RECT 547.890 4.690 548.270 5.070 ;
        RECT 548.550 4.690 548.930 5.070 ;
        RECT 549.590 4.690 549.970 5.070 ;
        RECT 550.590 4.690 550.970 5.070 ;
        RECT 551.250 4.690 551.630 5.070 ;
        RECT 551.910 4.690 552.290 5.070 ;
        RECT 552.830 4.690 553.210 5.070 ;
        RECT 553.490 4.690 553.870 5.070 ;
        RECT 554.150 4.690 554.530 5.070 ;
        RECT 555.070 4.690 555.450 5.070 ;
        RECT 555.730 4.690 556.110 5.070 ;
        RECT 556.390 4.690 556.770 5.070 ;
        RECT 557.310 4.690 557.690 5.070 ;
        RECT 557.970 4.690 558.350 5.070 ;
        RECT 558.630 4.690 559.010 5.070 ;
        RECT 559.550 4.690 559.930 5.070 ;
        RECT 560.210 4.690 560.590 5.070 ;
        RECT 560.870 4.690 561.250 5.070 ;
        RECT 561.790 4.690 562.170 5.070 ;
        RECT 562.450 4.690 562.830 5.070 ;
        RECT 563.110 4.690 563.490 5.070 ;
        RECT 564.030 4.690 564.410 5.070 ;
        RECT 564.690 4.690 565.070 5.070 ;
        RECT 565.350 4.690 565.730 5.070 ;
        RECT 566.370 4.690 566.750 5.070 ;
        RECT 567.030 4.690 567.410 5.070 ;
        RECT 567.690 4.690 568.070 5.070 ;
        RECT 569.750 4.690 570.130 5.070 ;
        RECT 570.750 4.690 571.130 5.070 ;
        RECT 571.410 4.690 571.790 5.070 ;
        RECT 572.070 4.690 572.450 5.070 ;
        RECT 572.990 4.690 573.370 5.070 ;
        RECT 573.650 4.690 574.030 5.070 ;
        RECT 574.310 4.690 574.690 5.070 ;
        RECT 575.230 4.690 575.610 5.070 ;
        RECT 575.890 4.690 576.270 5.070 ;
        RECT 576.550 4.690 576.930 5.070 ;
        RECT 577.470 4.690 577.850 5.070 ;
        RECT 578.130 4.690 578.510 5.070 ;
        RECT 578.790 4.690 579.170 5.070 ;
        RECT 579.710 4.690 580.090 5.070 ;
        RECT 580.370 4.690 580.750 5.070 ;
        RECT 581.030 4.690 581.410 5.070 ;
        RECT 581.950 4.690 582.330 5.070 ;
        RECT 582.610 4.690 582.990 5.070 ;
        RECT 583.270 4.690 583.650 5.070 ;
        RECT 584.190 4.690 584.570 5.070 ;
        RECT 584.850 4.690 585.230 5.070 ;
        RECT 585.510 4.690 585.890 5.070 ;
        RECT 586.430 4.690 586.810 5.070 ;
        RECT 587.090 4.690 587.470 5.070 ;
        RECT 587.750 4.690 588.130 5.070 ;
        RECT 588.670 4.690 589.050 5.070 ;
        RECT 589.330 4.690 589.710 5.070 ;
        RECT 589.990 4.690 590.370 5.070 ;
        RECT 591.030 4.690 591.410 5.070 ;
        RECT 592.030 4.690 592.410 5.070 ;
        RECT 592.690 4.690 593.070 5.070 ;
        RECT 593.350 4.690 593.730 5.070 ;
        RECT 594.270 4.690 594.650 5.070 ;
        RECT 594.930 4.690 595.310 5.070 ;
        RECT 595.590 4.690 595.970 5.070 ;
        RECT 596.510 4.690 596.890 5.070 ;
        RECT 597.170 4.690 597.550 5.070 ;
        RECT 597.830 4.690 598.210 5.070 ;
        RECT 598.750 4.690 599.130 5.070 ;
        RECT 599.410 4.690 599.790 5.070 ;
        RECT 600.070 4.690 600.450 5.070 ;
        RECT 600.990 4.690 601.370 5.070 ;
        RECT 601.650 4.690 602.030 5.070 ;
        RECT 602.310 4.690 602.690 5.070 ;
        RECT 603.230 4.690 603.610 5.070 ;
        RECT 603.890 4.690 604.270 5.070 ;
        RECT 604.550 4.690 604.930 5.070 ;
        RECT 605.470 4.690 605.850 5.070 ;
        RECT 606.130 4.690 606.510 5.070 ;
        RECT 606.790 4.690 607.170 5.070 ;
        RECT 607.810 4.690 608.190 5.070 ;
        RECT 608.470 4.690 608.850 5.070 ;
        RECT 609.130 4.690 609.510 5.070 ;
        RECT 611.190 4.690 611.570 5.070 ;
        RECT 612.190 4.690 612.570 5.070 ;
        RECT 612.850 4.690 613.230 5.070 ;
        RECT 613.510 4.690 613.890 5.070 ;
        RECT 614.430 4.690 614.810 5.070 ;
        RECT 615.090 4.690 615.470 5.070 ;
        RECT 615.750 4.690 616.130 5.070 ;
        RECT 616.670 4.690 617.050 5.070 ;
        RECT 617.330 4.690 617.710 5.070 ;
        RECT 617.990 4.690 618.370 5.070 ;
        RECT 618.910 4.690 619.290 5.070 ;
        RECT 619.570 4.690 619.950 5.070 ;
        RECT 620.230 4.690 620.610 5.070 ;
        RECT 621.150 4.690 621.530 5.070 ;
        RECT 621.810 4.690 622.190 5.070 ;
        RECT 622.470 4.690 622.850 5.070 ;
        RECT 623.390 4.690 623.770 5.070 ;
        RECT 624.050 4.690 624.430 5.070 ;
        RECT 624.710 4.690 625.090 5.070 ;
        RECT 625.630 4.690 626.010 5.070 ;
        RECT 626.290 4.690 626.670 5.070 ;
        RECT 626.950 4.690 627.330 5.070 ;
        RECT 627.870 4.690 628.250 5.070 ;
        RECT 628.530 4.690 628.910 5.070 ;
        RECT 629.190 4.690 629.570 5.070 ;
        RECT 630.110 4.690 630.490 5.070 ;
        RECT 630.770 4.690 631.150 5.070 ;
        RECT 631.430 4.690 631.810 5.070 ;
        RECT 632.470 4.690 632.850 5.070 ;
        RECT 633.470 4.690 633.850 5.070 ;
        RECT 634.130 4.690 634.510 5.070 ;
        RECT 634.790 4.690 635.170 5.070 ;
        RECT 635.710 4.690 636.090 5.070 ;
        RECT 636.370 4.690 636.750 5.070 ;
        RECT 637.030 4.690 637.410 5.070 ;
        RECT 637.950 4.690 638.330 5.070 ;
        RECT 638.610 4.690 638.990 5.070 ;
        RECT 639.270 4.690 639.650 5.070 ;
        RECT 640.190 4.690 640.570 5.070 ;
        RECT 640.850 4.690 641.230 5.070 ;
        RECT 641.510 4.690 641.890 5.070 ;
        RECT 642.430 4.690 642.810 5.070 ;
        RECT 643.090 4.690 643.470 5.070 ;
        RECT 643.750 4.690 644.130 5.070 ;
        RECT 644.670 4.690 645.050 5.070 ;
        RECT 645.330 4.690 645.710 5.070 ;
        RECT 645.990 4.690 646.370 5.070 ;
        RECT 646.910 4.690 647.290 5.070 ;
        RECT 647.570 4.690 647.950 5.070 ;
        RECT 648.230 4.690 648.610 5.070 ;
        RECT 649.150 4.690 649.530 5.070 ;
        RECT 649.810 4.690 650.190 5.070 ;
        RECT 650.470 4.690 650.850 5.070 ;
        RECT 651.490 4.690 651.870 5.070 ;
        RECT 652.150 4.690 652.530 5.070 ;
        RECT 652.810 4.690 653.190 5.070 ;
        RECT 654.870 4.690 655.250 5.070 ;
        RECT 655.870 4.690 656.250 5.070 ;
        RECT 656.530 4.690 656.910 5.070 ;
        RECT 657.190 4.690 657.570 5.070 ;
        RECT 658.110 4.690 658.490 5.070 ;
        RECT 658.770 4.690 659.150 5.070 ;
        RECT 659.430 4.690 659.810 5.070 ;
        RECT 660.350 4.690 660.730 5.070 ;
        RECT 661.010 4.690 661.390 5.070 ;
        RECT 661.670 4.690 662.050 5.070 ;
        RECT 662.590 4.690 662.970 5.070 ;
        RECT 663.250 4.690 663.630 5.070 ;
        RECT 663.910 4.690 664.290 5.070 ;
        RECT 664.830 4.690 665.210 5.070 ;
        RECT 665.490 4.690 665.870 5.070 ;
        RECT 666.150 4.690 666.530 5.070 ;
        RECT 667.070 4.690 667.450 5.070 ;
        RECT 667.730 4.690 668.110 5.070 ;
        RECT 668.390 4.690 668.770 5.070 ;
        RECT 669.310 4.690 669.690 5.070 ;
        RECT 669.970 4.690 670.350 5.070 ;
        RECT 670.630 4.690 671.010 5.070 ;
        RECT 671.550 4.690 671.930 5.070 ;
        RECT 672.210 4.690 672.590 5.070 ;
        RECT 672.870 4.690 673.250 5.070 ;
        RECT 673.790 4.690 674.170 5.070 ;
        RECT 674.450 4.690 674.830 5.070 ;
        RECT 675.110 4.690 675.490 5.070 ;
        RECT 676.150 4.690 676.530 5.070 ;
        RECT 677.150 4.690 677.530 5.070 ;
        RECT 677.810 4.690 678.190 5.070 ;
        RECT 678.470 4.690 678.850 5.070 ;
        RECT 679.490 4.690 679.870 5.070 ;
        RECT 0.850 0.770 1.230 1.150 ;
        RECT 1.990 0.770 2.370 1.150 ;
        RECT 7.430 0.770 7.810 1.150 ;
        RECT 8.090 0.770 8.470 1.150 ;
        RECT 8.750 0.770 9.130 1.150 ;
        RECT 14.300 0.770 14.680 1.150 ;
        RECT 15.620 0.770 16.000 1.150 ;
        RECT 17.660 0.770 18.040 1.150 ;
        RECT 18.980 0.770 19.360 1.150 ;
        RECT 25.620 0.770 26.000 1.150 ;
        RECT 26.280 0.770 26.660 1.150 ;
        RECT 26.940 0.770 27.320 1.150 ;
        RECT 32.490 0.770 32.870 1.150 ;
        RECT 33.810 0.770 34.190 1.150 ;
        RECT 36.130 0.770 36.510 1.150 ;
        RECT 41.570 0.770 41.950 1.150 ;
        RECT 42.230 0.770 42.610 1.150 ;
        RECT 42.890 0.770 43.270 1.150 ;
        RECT 48.440 0.770 48.820 1.150 ;
        RECT 49.760 0.770 50.140 1.150 ;
        RECT 56.400 0.770 56.780 1.150 ;
        RECT 57.060 0.770 57.440 1.150 ;
        RECT 57.720 0.770 58.100 1.150 ;
        RECT 63.270 0.770 63.650 1.150 ;
        RECT 64.590 0.770 64.970 1.150 ;
        RECT 66.630 0.770 67.010 1.150 ;
        RECT 67.950 0.770 68.330 1.150 ;
        RECT 70.270 0.770 70.650 1.150 ;
        RECT 75.710 0.770 76.090 1.150 ;
        RECT 76.370 0.770 76.750 1.150 ;
        RECT 77.030 0.770 77.410 1.150 ;
        RECT 82.580 0.770 82.960 1.150 ;
        RECT 83.900 0.770 84.280 1.150 ;
        RECT 90.540 0.770 90.920 1.150 ;
        RECT 91.200 0.770 91.580 1.150 ;
        RECT 91.860 0.770 92.240 1.150 ;
        RECT 97.410 0.770 97.790 1.150 ;
        RECT 98.730 0.770 99.110 1.150 ;
        RECT 100.770 0.770 101.150 1.150 ;
        RECT 102.090 0.770 102.470 1.150 ;
        RECT 104.410 0.770 104.790 1.150 ;
        RECT 109.850 0.770 110.230 1.150 ;
        RECT 110.510 0.770 110.890 1.150 ;
        RECT 111.170 0.770 111.550 1.150 ;
        RECT 116.720 0.770 117.100 1.150 ;
        RECT 118.040 0.770 118.420 1.150 ;
        RECT 124.680 0.770 125.060 1.150 ;
        RECT 125.340 0.770 125.720 1.150 ;
        RECT 126.000 0.770 126.380 1.150 ;
        RECT 131.550 0.770 131.930 1.150 ;
        RECT 132.870 0.770 133.250 1.150 ;
        RECT 135.190 0.770 135.570 1.150 ;
        RECT 136.190 0.770 136.570 1.150 ;
        RECT 136.850 0.770 137.230 1.150 ;
        RECT 137.510 0.770 137.890 1.150 ;
        RECT 138.430 0.770 138.810 1.150 ;
        RECT 139.090 0.770 139.470 1.150 ;
        RECT 139.750 0.770 140.130 1.150 ;
        RECT 140.510 0.770 140.890 1.150 ;
        RECT 141.830 0.770 142.210 1.150 ;
        RECT 144.030 0.770 144.410 1.150 ;
        RECT 144.690 0.770 145.070 1.150 ;
        RECT 145.350 0.770 145.730 1.150 ;
        RECT 146.270 0.770 146.650 1.150 ;
        RECT 146.930 0.770 147.310 1.150 ;
        RECT 147.590 0.770 147.970 1.150 ;
        RECT 148.510 0.770 148.890 1.150 ;
        RECT 149.170 0.770 149.550 1.150 ;
        RECT 149.830 0.770 150.210 1.150 ;
        RECT 150.750 0.770 151.130 1.150 ;
        RECT 151.410 0.770 151.790 1.150 ;
        RECT 152.070 0.770 152.450 1.150 ;
        RECT 152.990 0.770 153.370 1.150 ;
        RECT 153.650 0.770 154.030 1.150 ;
        RECT 154.310 0.770 154.690 1.150 ;
        RECT 155.350 0.770 155.730 1.150 ;
        RECT 156.350 0.770 156.730 1.150 ;
        RECT 157.010 0.770 157.390 1.150 ;
        RECT 157.670 0.770 158.050 1.150 ;
        RECT 158.590 0.770 158.970 1.150 ;
        RECT 159.250 0.770 159.630 1.150 ;
        RECT 159.910 0.770 160.290 1.150 ;
        RECT 160.830 0.770 161.210 1.150 ;
        RECT 161.490 0.770 161.870 1.150 ;
        RECT 162.150 0.770 162.530 1.150 ;
        RECT 163.070 0.770 163.450 1.150 ;
        RECT 163.730 0.770 164.110 1.150 ;
        RECT 164.390 0.770 164.770 1.150 ;
        RECT 165.310 0.770 165.690 1.150 ;
        RECT 165.970 0.770 166.350 1.150 ;
        RECT 166.630 0.770 167.010 1.150 ;
        RECT 167.550 0.770 167.930 1.150 ;
        RECT 168.210 0.770 168.590 1.150 ;
        RECT 168.870 0.770 169.250 1.150 ;
        RECT 169.790 0.770 170.170 1.150 ;
        RECT 170.450 0.770 170.830 1.150 ;
        RECT 171.110 0.770 171.490 1.150 ;
        RECT 172.030 0.770 172.410 1.150 ;
        RECT 172.690 0.770 173.070 1.150 ;
        RECT 173.350 0.770 173.730 1.150 ;
        RECT 174.270 0.770 174.650 1.150 ;
        RECT 174.930 0.770 175.310 1.150 ;
        RECT 175.590 0.770 175.970 1.150 ;
        RECT 176.630 0.770 177.010 1.150 ;
        RECT 177.630 0.770 178.010 1.150 ;
        RECT 178.290 0.770 178.670 1.150 ;
        RECT 178.950 0.770 179.330 1.150 ;
        RECT 179.870 0.770 180.250 1.150 ;
        RECT 180.530 0.770 180.910 1.150 ;
        RECT 181.190 0.770 181.570 1.150 ;
        RECT 181.950 0.770 182.330 1.150 ;
        RECT 183.270 0.770 183.650 1.150 ;
        RECT 185.470 0.770 185.850 1.150 ;
        RECT 186.130 0.770 186.510 1.150 ;
        RECT 186.790 0.770 187.170 1.150 ;
        RECT 187.710 0.770 188.090 1.150 ;
        RECT 188.370 0.770 188.750 1.150 ;
        RECT 189.030 0.770 189.410 1.150 ;
        RECT 189.950 0.770 190.330 1.150 ;
        RECT 190.610 0.770 190.990 1.150 ;
        RECT 191.270 0.770 191.650 1.150 ;
        RECT 192.190 0.770 192.570 1.150 ;
        RECT 192.850 0.770 193.230 1.150 ;
        RECT 193.510 0.770 193.890 1.150 ;
        RECT 194.430 0.770 194.810 1.150 ;
        RECT 195.090 0.770 195.470 1.150 ;
        RECT 195.750 0.770 196.130 1.150 ;
        RECT 196.790 0.770 197.170 1.150 ;
        RECT 197.790 0.770 198.170 1.150 ;
        RECT 198.450 0.770 198.830 1.150 ;
        RECT 199.110 0.770 199.490 1.150 ;
        RECT 200.030 0.770 200.410 1.150 ;
        RECT 200.690 0.770 201.070 1.150 ;
        RECT 201.350 0.770 201.730 1.150 ;
        RECT 202.270 0.770 202.650 1.150 ;
        RECT 202.930 0.770 203.310 1.150 ;
        RECT 203.590 0.770 203.970 1.150 ;
        RECT 204.510 0.770 204.890 1.150 ;
        RECT 205.170 0.770 205.550 1.150 ;
        RECT 205.830 0.770 206.210 1.150 ;
        RECT 206.750 0.770 207.130 1.150 ;
        RECT 207.410 0.770 207.790 1.150 ;
        RECT 208.070 0.770 208.450 1.150 ;
        RECT 208.990 0.770 209.370 1.150 ;
        RECT 209.650 0.770 210.030 1.150 ;
        RECT 210.310 0.770 210.690 1.150 ;
        RECT 211.230 0.770 211.610 1.150 ;
        RECT 211.890 0.770 212.270 1.150 ;
        RECT 212.550 0.770 212.930 1.150 ;
        RECT 213.470 0.770 213.850 1.150 ;
        RECT 214.130 0.770 214.510 1.150 ;
        RECT 214.790 0.770 215.170 1.150 ;
        RECT 215.710 0.770 216.090 1.150 ;
        RECT 216.370 0.770 216.750 1.150 ;
        RECT 217.030 0.770 217.410 1.150 ;
        RECT 218.070 0.770 218.450 1.150 ;
        RECT 219.070 0.770 219.450 1.150 ;
        RECT 219.730 0.770 220.110 1.150 ;
        RECT 220.390 0.770 220.770 1.150 ;
        RECT 221.310 0.770 221.690 1.150 ;
        RECT 221.970 0.770 222.350 1.150 ;
        RECT 222.630 0.770 223.010 1.150 ;
        RECT 223.550 0.770 223.930 1.150 ;
        RECT 224.210 0.770 224.590 1.150 ;
        RECT 224.870 0.770 225.250 1.150 ;
        RECT 225.630 0.770 226.010 1.150 ;
        RECT 226.950 0.770 227.330 1.150 ;
        RECT 229.150 0.770 229.530 1.150 ;
        RECT 229.810 0.770 230.190 1.150 ;
        RECT 230.470 0.770 230.850 1.150 ;
        RECT 231.390 0.770 231.770 1.150 ;
        RECT 232.050 0.770 232.430 1.150 ;
        RECT 232.710 0.770 233.090 1.150 ;
        RECT 233.630 0.770 234.010 1.150 ;
        RECT 234.290 0.770 234.670 1.150 ;
        RECT 234.950 0.770 235.330 1.150 ;
        RECT 235.870 0.770 236.250 1.150 ;
        RECT 236.530 0.770 236.910 1.150 ;
        RECT 237.190 0.770 237.570 1.150 ;
        RECT 238.230 0.770 238.610 1.150 ;
        RECT 239.230 0.770 239.610 1.150 ;
        RECT 239.890 0.770 240.270 1.150 ;
        RECT 240.550 0.770 240.930 1.150 ;
        RECT 241.470 0.770 241.850 1.150 ;
        RECT 242.130 0.770 242.510 1.150 ;
        RECT 242.790 0.770 243.170 1.150 ;
        RECT 243.710 0.770 244.090 1.150 ;
        RECT 244.370 0.770 244.750 1.150 ;
        RECT 245.030 0.770 245.410 1.150 ;
        RECT 245.950 0.770 246.330 1.150 ;
        RECT 246.610 0.770 246.990 1.150 ;
        RECT 247.270 0.770 247.650 1.150 ;
        RECT 248.190 0.770 248.570 1.150 ;
        RECT 248.850 0.770 249.230 1.150 ;
        RECT 249.510 0.770 249.890 1.150 ;
        RECT 250.430 0.770 250.810 1.150 ;
        RECT 251.090 0.770 251.470 1.150 ;
        RECT 251.750 0.770 252.130 1.150 ;
        RECT 252.670 0.770 253.050 1.150 ;
        RECT 253.330 0.770 253.710 1.150 ;
        RECT 253.990 0.770 254.370 1.150 ;
        RECT 254.910 0.770 255.290 1.150 ;
        RECT 255.570 0.770 255.950 1.150 ;
        RECT 256.230 0.770 256.610 1.150 ;
        RECT 257.150 0.770 257.530 1.150 ;
        RECT 257.810 0.770 258.190 1.150 ;
        RECT 258.470 0.770 258.850 1.150 ;
        RECT 259.510 0.770 259.890 1.150 ;
        RECT 260.510 0.770 260.890 1.150 ;
        RECT 261.170 0.770 261.550 1.150 ;
        RECT 261.830 0.770 262.210 1.150 ;
        RECT 262.750 0.770 263.130 1.150 ;
        RECT 263.410 0.770 263.790 1.150 ;
        RECT 264.070 0.770 264.450 1.150 ;
        RECT 264.990 0.770 265.370 1.150 ;
        RECT 265.650 0.770 266.030 1.150 ;
        RECT 266.310 0.770 266.690 1.150 ;
        RECT 267.070 0.770 267.450 1.150 ;
        RECT 268.390 0.770 268.770 1.150 ;
        RECT 270.590 0.770 270.970 1.150 ;
        RECT 271.250 0.770 271.630 1.150 ;
        RECT 271.910 0.770 272.290 1.150 ;
        RECT 272.830 0.770 273.210 1.150 ;
        RECT 273.490 0.770 273.870 1.150 ;
        RECT 274.150 0.770 274.530 1.150 ;
        RECT 275.070 0.770 275.450 1.150 ;
        RECT 275.730 0.770 276.110 1.150 ;
        RECT 276.390 0.770 276.770 1.150 ;
        RECT 277.310 0.770 277.690 1.150 ;
        RECT 277.970 0.770 278.350 1.150 ;
        RECT 278.630 0.770 279.010 1.150 ;
        RECT 279.670 0.770 280.050 1.150 ;
        RECT 280.670 0.770 281.050 1.150 ;
        RECT 281.330 0.770 281.710 1.150 ;
        RECT 281.990 0.770 282.370 1.150 ;
        RECT 282.910 0.770 283.290 1.150 ;
        RECT 283.570 0.770 283.950 1.150 ;
        RECT 284.230 0.770 284.610 1.150 ;
        RECT 285.150 0.770 285.530 1.150 ;
        RECT 285.810 0.770 286.190 1.150 ;
        RECT 286.470 0.770 286.850 1.150 ;
        RECT 287.390 0.770 287.770 1.150 ;
        RECT 288.050 0.770 288.430 1.150 ;
        RECT 288.710 0.770 289.090 1.150 ;
        RECT 289.630 0.770 290.010 1.150 ;
        RECT 290.290 0.770 290.670 1.150 ;
        RECT 290.950 0.770 291.330 1.150 ;
        RECT 291.870 0.770 292.250 1.150 ;
        RECT 292.530 0.770 292.910 1.150 ;
        RECT 293.190 0.770 293.570 1.150 ;
        RECT 294.110 0.770 294.490 1.150 ;
        RECT 294.770 0.770 295.150 1.150 ;
        RECT 295.430 0.770 295.810 1.150 ;
        RECT 296.350 0.770 296.730 1.150 ;
        RECT 297.010 0.770 297.390 1.150 ;
        RECT 297.670 0.770 298.050 1.150 ;
        RECT 298.590 0.770 298.970 1.150 ;
        RECT 299.250 0.770 299.630 1.150 ;
        RECT 299.910 0.770 300.290 1.150 ;
        RECT 300.950 0.770 301.330 1.150 ;
        RECT 301.950 0.770 302.330 1.150 ;
        RECT 302.610 0.770 302.990 1.150 ;
        RECT 303.270 0.770 303.650 1.150 ;
        RECT 304.190 0.770 304.570 1.150 ;
        RECT 304.850 0.770 305.230 1.150 ;
        RECT 305.510 0.770 305.890 1.150 ;
        RECT 306.430 0.770 306.810 1.150 ;
        RECT 307.090 0.770 307.470 1.150 ;
        RECT 307.750 0.770 308.130 1.150 ;
        RECT 308.670 0.770 309.050 1.150 ;
        RECT 309.330 0.770 309.710 1.150 ;
        RECT 309.990 0.770 310.370 1.150 ;
        RECT 310.750 0.770 311.130 1.150 ;
        RECT 312.070 0.770 312.450 1.150 ;
        RECT 314.270 0.770 314.650 1.150 ;
        RECT 314.930 0.770 315.310 1.150 ;
        RECT 315.590 0.770 315.970 1.150 ;
        RECT 316.510 0.770 316.890 1.150 ;
        RECT 317.170 0.770 317.550 1.150 ;
        RECT 317.830 0.770 318.210 1.150 ;
        RECT 318.750 0.770 319.130 1.150 ;
        RECT 319.410 0.770 319.790 1.150 ;
        RECT 320.070 0.770 320.450 1.150 ;
        RECT 321.110 0.770 321.490 1.150 ;
        RECT 322.110 0.770 322.490 1.150 ;
        RECT 322.770 0.770 323.150 1.150 ;
        RECT 323.430 0.770 323.810 1.150 ;
        RECT 324.350 0.770 324.730 1.150 ;
        RECT 325.010 0.770 325.390 1.150 ;
        RECT 325.670 0.770 326.050 1.150 ;
        RECT 326.590 0.770 326.970 1.150 ;
        RECT 327.250 0.770 327.630 1.150 ;
        RECT 327.910 0.770 328.290 1.150 ;
        RECT 328.830 0.770 329.210 1.150 ;
        RECT 329.490 0.770 329.870 1.150 ;
        RECT 330.150 0.770 330.530 1.150 ;
        RECT 331.070 0.770 331.450 1.150 ;
        RECT 331.730 0.770 332.110 1.150 ;
        RECT 332.390 0.770 332.770 1.150 ;
        RECT 333.310 0.770 333.690 1.150 ;
        RECT 333.970 0.770 334.350 1.150 ;
        RECT 334.630 0.770 335.010 1.150 ;
        RECT 335.550 0.770 335.930 1.150 ;
        RECT 336.210 0.770 336.590 1.150 ;
        RECT 336.870 0.770 337.250 1.150 ;
        RECT 337.790 0.770 338.170 1.150 ;
        RECT 338.450 0.770 338.830 1.150 ;
        RECT 339.110 0.770 339.490 1.150 ;
        RECT 340.030 0.770 340.410 1.150 ;
        RECT 340.690 0.770 341.070 1.150 ;
        RECT 341.350 0.770 341.730 1.150 ;
        RECT 342.390 0.770 342.770 1.150 ;
        RECT 343.390 0.770 343.770 1.150 ;
        RECT 344.050 0.770 344.430 1.150 ;
        RECT 344.710 0.770 345.090 1.150 ;
        RECT 345.630 0.770 346.010 1.150 ;
        RECT 346.290 0.770 346.670 1.150 ;
        RECT 346.950 0.770 347.330 1.150 ;
        RECT 347.870 0.770 348.250 1.150 ;
        RECT 348.530 0.770 348.910 1.150 ;
        RECT 349.190 0.770 349.570 1.150 ;
        RECT 350.110 0.770 350.490 1.150 ;
        RECT 350.770 0.770 351.150 1.150 ;
        RECT 351.430 0.770 351.810 1.150 ;
        RECT 352.190 0.770 352.570 1.150 ;
        RECT 353.510 0.770 353.890 1.150 ;
        RECT 355.710 0.770 356.090 1.150 ;
        RECT 356.370 0.770 356.750 1.150 ;
        RECT 357.030 0.770 357.410 1.150 ;
        RECT 357.950 0.770 358.330 1.150 ;
        RECT 358.610 0.770 358.990 1.150 ;
        RECT 359.270 0.770 359.650 1.150 ;
        RECT 360.190 0.770 360.570 1.150 ;
        RECT 360.850 0.770 361.230 1.150 ;
        RECT 361.510 0.770 361.890 1.150 ;
        RECT 362.550 0.770 362.930 1.150 ;
        RECT 363.550 0.770 363.930 1.150 ;
        RECT 364.210 0.770 364.590 1.150 ;
        RECT 364.870 0.770 365.250 1.150 ;
        RECT 365.790 0.770 366.170 1.150 ;
        RECT 366.450 0.770 366.830 1.150 ;
        RECT 367.110 0.770 367.490 1.150 ;
        RECT 368.030 0.770 368.410 1.150 ;
        RECT 368.690 0.770 369.070 1.150 ;
        RECT 369.350 0.770 369.730 1.150 ;
        RECT 370.270 0.770 370.650 1.150 ;
        RECT 370.930 0.770 371.310 1.150 ;
        RECT 371.590 0.770 371.970 1.150 ;
        RECT 372.510 0.770 372.890 1.150 ;
        RECT 373.170 0.770 373.550 1.150 ;
        RECT 373.830 0.770 374.210 1.150 ;
        RECT 374.750 0.770 375.130 1.150 ;
        RECT 375.410 0.770 375.790 1.150 ;
        RECT 376.070 0.770 376.450 1.150 ;
        RECT 376.990 0.770 377.370 1.150 ;
        RECT 377.650 0.770 378.030 1.150 ;
        RECT 378.310 0.770 378.690 1.150 ;
        RECT 379.230 0.770 379.610 1.150 ;
        RECT 379.890 0.770 380.270 1.150 ;
        RECT 380.550 0.770 380.930 1.150 ;
        RECT 381.470 0.770 381.850 1.150 ;
        RECT 382.130 0.770 382.510 1.150 ;
        RECT 382.790 0.770 383.170 1.150 ;
        RECT 383.830 0.770 384.210 1.150 ;
        RECT 384.830 0.770 385.210 1.150 ;
        RECT 385.490 0.770 385.870 1.150 ;
        RECT 386.150 0.770 386.530 1.150 ;
        RECT 387.070 0.770 387.450 1.150 ;
        RECT 387.730 0.770 388.110 1.150 ;
        RECT 388.390 0.770 388.770 1.150 ;
        RECT 389.310 0.770 389.690 1.150 ;
        RECT 389.970 0.770 390.350 1.150 ;
        RECT 390.630 0.770 391.010 1.150 ;
        RECT 391.550 0.770 391.930 1.150 ;
        RECT 392.210 0.770 392.590 1.150 ;
        RECT 392.870 0.770 393.250 1.150 ;
        RECT 393.790 0.770 394.170 1.150 ;
        RECT 394.450 0.770 394.830 1.150 ;
        RECT 395.110 0.770 395.490 1.150 ;
        RECT 395.870 0.770 396.250 1.150 ;
        RECT 397.190 0.770 397.570 1.150 ;
        RECT 399.390 0.770 399.770 1.150 ;
        RECT 400.050 0.770 400.430 1.150 ;
        RECT 400.710 0.770 401.090 1.150 ;
        RECT 401.630 0.770 402.010 1.150 ;
        RECT 402.290 0.770 402.670 1.150 ;
        RECT 402.950 0.770 403.330 1.150 ;
        RECT 403.990 0.770 404.370 1.150 ;
        RECT 404.990 0.770 405.370 1.150 ;
        RECT 405.650 0.770 406.030 1.150 ;
        RECT 406.310 0.770 406.690 1.150 ;
        RECT 407.230 0.770 407.610 1.150 ;
        RECT 407.890 0.770 408.270 1.150 ;
        RECT 408.550 0.770 408.930 1.150 ;
        RECT 409.470 0.770 409.850 1.150 ;
        RECT 410.130 0.770 410.510 1.150 ;
        RECT 410.790 0.770 411.170 1.150 ;
        RECT 411.710 0.770 412.090 1.150 ;
        RECT 412.370 0.770 412.750 1.150 ;
        RECT 413.030 0.770 413.410 1.150 ;
        RECT 413.950 0.770 414.330 1.150 ;
        RECT 414.610 0.770 414.990 1.150 ;
        RECT 415.270 0.770 415.650 1.150 ;
        RECT 416.190 0.770 416.570 1.150 ;
        RECT 416.850 0.770 417.230 1.150 ;
        RECT 417.510 0.770 417.890 1.150 ;
        RECT 418.430 0.770 418.810 1.150 ;
        RECT 419.090 0.770 419.470 1.150 ;
        RECT 419.750 0.770 420.130 1.150 ;
        RECT 420.670 0.770 421.050 1.150 ;
        RECT 421.330 0.770 421.710 1.150 ;
        RECT 421.990 0.770 422.370 1.150 ;
        RECT 422.910 0.770 423.290 1.150 ;
        RECT 423.570 0.770 423.950 1.150 ;
        RECT 424.230 0.770 424.610 1.150 ;
        RECT 425.270 0.770 425.650 1.150 ;
        RECT 426.270 0.770 426.650 1.150 ;
        RECT 426.930 0.770 427.310 1.150 ;
        RECT 427.590 0.770 427.970 1.150 ;
        RECT 428.510 0.770 428.890 1.150 ;
        RECT 429.170 0.770 429.550 1.150 ;
        RECT 429.830 0.770 430.210 1.150 ;
        RECT 430.750 0.770 431.130 1.150 ;
        RECT 431.410 0.770 431.790 1.150 ;
        RECT 432.070 0.770 432.450 1.150 ;
        RECT 432.990 0.770 433.370 1.150 ;
        RECT 433.650 0.770 434.030 1.150 ;
        RECT 434.310 0.770 434.690 1.150 ;
        RECT 435.230 0.770 435.610 1.150 ;
        RECT 435.890 0.770 436.270 1.150 ;
        RECT 436.550 0.770 436.930 1.150 ;
        RECT 437.310 0.770 437.690 1.150 ;
        RECT 438.630 0.770 439.010 1.150 ;
        RECT 440.830 0.770 441.210 1.150 ;
        RECT 441.490 0.770 441.870 1.150 ;
        RECT 442.150 0.770 442.530 1.150 ;
        RECT 443.070 0.770 443.450 1.150 ;
        RECT 443.730 0.770 444.110 1.150 ;
        RECT 444.390 0.770 444.770 1.150 ;
        RECT 445.430 0.770 445.810 1.150 ;
        RECT 446.430 0.770 446.810 1.150 ;
        RECT 447.090 0.770 447.470 1.150 ;
        RECT 447.750 0.770 448.130 1.150 ;
        RECT 448.670 0.770 449.050 1.150 ;
        RECT 449.330 0.770 449.710 1.150 ;
        RECT 449.990 0.770 450.370 1.150 ;
        RECT 450.910 0.770 451.290 1.150 ;
        RECT 451.570 0.770 451.950 1.150 ;
        RECT 452.230 0.770 452.610 1.150 ;
        RECT 453.150 0.770 453.530 1.150 ;
        RECT 453.810 0.770 454.190 1.150 ;
        RECT 454.470 0.770 454.850 1.150 ;
        RECT 455.390 0.770 455.770 1.150 ;
        RECT 456.050 0.770 456.430 1.150 ;
        RECT 456.710 0.770 457.090 1.150 ;
        RECT 457.630 0.770 458.010 1.150 ;
        RECT 458.290 0.770 458.670 1.150 ;
        RECT 458.950 0.770 459.330 1.150 ;
        RECT 459.870 0.770 460.250 1.150 ;
        RECT 460.530 0.770 460.910 1.150 ;
        RECT 461.190 0.770 461.570 1.150 ;
        RECT 462.110 0.770 462.490 1.150 ;
        RECT 462.770 0.770 463.150 1.150 ;
        RECT 463.430 0.770 463.810 1.150 ;
        RECT 464.350 0.770 464.730 1.150 ;
        RECT 465.010 0.770 465.390 1.150 ;
        RECT 465.670 0.770 466.050 1.150 ;
        RECT 466.710 0.770 467.090 1.150 ;
        RECT 467.710 0.770 468.090 1.150 ;
        RECT 468.370 0.770 468.750 1.150 ;
        RECT 469.030 0.770 469.410 1.150 ;
        RECT 469.950 0.770 470.330 1.150 ;
        RECT 470.610 0.770 470.990 1.150 ;
        RECT 471.270 0.770 471.650 1.150 ;
        RECT 472.190 0.770 472.570 1.150 ;
        RECT 472.850 0.770 473.230 1.150 ;
        RECT 473.510 0.770 473.890 1.150 ;
        RECT 474.430 0.770 474.810 1.150 ;
        RECT 475.090 0.770 475.470 1.150 ;
        RECT 475.750 0.770 476.130 1.150 ;
        RECT 476.670 0.770 477.050 1.150 ;
        RECT 477.330 0.770 477.710 1.150 ;
        RECT 477.990 0.770 478.370 1.150 ;
        RECT 478.910 0.770 479.290 1.150 ;
        RECT 479.570 0.770 479.950 1.150 ;
        RECT 480.230 0.770 480.610 1.150 ;
        RECT 480.990 0.770 481.370 1.150 ;
        RECT 482.310 0.770 482.690 1.150 ;
        RECT 484.510 0.770 484.890 1.150 ;
        RECT 485.170 0.770 485.550 1.150 ;
        RECT 485.830 0.770 486.210 1.150 ;
        RECT 486.870 0.770 487.250 1.150 ;
        RECT 487.870 0.770 488.250 1.150 ;
        RECT 488.530 0.770 488.910 1.150 ;
        RECT 489.190 0.770 489.570 1.150 ;
        RECT 490.110 0.770 490.490 1.150 ;
        RECT 490.770 0.770 491.150 1.150 ;
        RECT 491.430 0.770 491.810 1.150 ;
        RECT 492.350 0.770 492.730 1.150 ;
        RECT 493.010 0.770 493.390 1.150 ;
        RECT 493.670 0.770 494.050 1.150 ;
        RECT 494.590 0.770 494.970 1.150 ;
        RECT 495.250 0.770 495.630 1.150 ;
        RECT 495.910 0.770 496.290 1.150 ;
        RECT 496.830 0.770 497.210 1.150 ;
        RECT 497.490 0.770 497.870 1.150 ;
        RECT 498.150 0.770 498.530 1.150 ;
        RECT 499.070 0.770 499.450 1.150 ;
        RECT 499.730 0.770 500.110 1.150 ;
        RECT 500.390 0.770 500.770 1.150 ;
        RECT 501.310 0.770 501.690 1.150 ;
        RECT 501.970 0.770 502.350 1.150 ;
        RECT 502.630 0.770 503.010 1.150 ;
        RECT 503.550 0.770 503.930 1.150 ;
        RECT 504.210 0.770 504.590 1.150 ;
        RECT 504.870 0.770 505.250 1.150 ;
        RECT 505.790 0.770 506.170 1.150 ;
        RECT 506.450 0.770 506.830 1.150 ;
        RECT 507.110 0.770 507.490 1.150 ;
        RECT 508.150 0.770 508.530 1.150 ;
        RECT 509.150 0.770 509.530 1.150 ;
        RECT 509.810 0.770 510.190 1.150 ;
        RECT 510.470 0.770 510.850 1.150 ;
        RECT 511.390 0.770 511.770 1.150 ;
        RECT 512.050 0.770 512.430 1.150 ;
        RECT 512.710 0.770 513.090 1.150 ;
        RECT 513.630 0.770 514.010 1.150 ;
        RECT 514.290 0.770 514.670 1.150 ;
        RECT 514.950 0.770 515.330 1.150 ;
        RECT 515.870 0.770 516.250 1.150 ;
        RECT 516.530 0.770 516.910 1.150 ;
        RECT 517.190 0.770 517.570 1.150 ;
        RECT 518.110 0.770 518.490 1.150 ;
        RECT 518.770 0.770 519.150 1.150 ;
        RECT 519.430 0.770 519.810 1.150 ;
        RECT 520.350 0.770 520.730 1.150 ;
        RECT 521.010 0.770 521.390 1.150 ;
        RECT 521.670 0.770 522.050 1.150 ;
        RECT 522.430 0.770 522.810 1.150 ;
        RECT 523.750 0.770 524.130 1.150 ;
        RECT 525.950 0.770 526.330 1.150 ;
        RECT 526.610 0.770 526.990 1.150 ;
        RECT 527.270 0.770 527.650 1.150 ;
        RECT 528.310 0.770 528.690 1.150 ;
        RECT 529.310 0.770 529.690 1.150 ;
        RECT 529.970 0.770 530.350 1.150 ;
        RECT 530.630 0.770 531.010 1.150 ;
        RECT 531.550 0.770 531.930 1.150 ;
        RECT 532.210 0.770 532.590 1.150 ;
        RECT 532.870 0.770 533.250 1.150 ;
        RECT 533.790 0.770 534.170 1.150 ;
        RECT 534.450 0.770 534.830 1.150 ;
        RECT 535.110 0.770 535.490 1.150 ;
        RECT 536.030 0.770 536.410 1.150 ;
        RECT 536.690 0.770 537.070 1.150 ;
        RECT 537.350 0.770 537.730 1.150 ;
        RECT 538.270 0.770 538.650 1.150 ;
        RECT 538.930 0.770 539.310 1.150 ;
        RECT 539.590 0.770 539.970 1.150 ;
        RECT 540.510 0.770 540.890 1.150 ;
        RECT 541.170 0.770 541.550 1.150 ;
        RECT 541.830 0.770 542.210 1.150 ;
        RECT 542.750 0.770 543.130 1.150 ;
        RECT 543.410 0.770 543.790 1.150 ;
        RECT 544.070 0.770 544.450 1.150 ;
        RECT 544.990 0.770 545.370 1.150 ;
        RECT 545.650 0.770 546.030 1.150 ;
        RECT 546.310 0.770 546.690 1.150 ;
        RECT 547.230 0.770 547.610 1.150 ;
        RECT 547.890 0.770 548.270 1.150 ;
        RECT 548.550 0.770 548.930 1.150 ;
        RECT 549.590 0.770 549.970 1.150 ;
        RECT 550.590 0.770 550.970 1.150 ;
        RECT 551.250 0.770 551.630 1.150 ;
        RECT 551.910 0.770 552.290 1.150 ;
        RECT 552.830 0.770 553.210 1.150 ;
        RECT 553.490 0.770 553.870 1.150 ;
        RECT 554.150 0.770 554.530 1.150 ;
        RECT 555.070 0.770 555.450 1.150 ;
        RECT 555.730 0.770 556.110 1.150 ;
        RECT 556.390 0.770 556.770 1.150 ;
        RECT 557.310 0.770 557.690 1.150 ;
        RECT 557.970 0.770 558.350 1.150 ;
        RECT 558.630 0.770 559.010 1.150 ;
        RECT 559.550 0.770 559.930 1.150 ;
        RECT 560.210 0.770 560.590 1.150 ;
        RECT 560.870 0.770 561.250 1.150 ;
        RECT 561.790 0.770 562.170 1.150 ;
        RECT 562.450 0.770 562.830 1.150 ;
        RECT 563.110 0.770 563.490 1.150 ;
        RECT 564.030 0.770 564.410 1.150 ;
        RECT 564.690 0.770 565.070 1.150 ;
        RECT 565.350 0.770 565.730 1.150 ;
        RECT 566.110 0.770 566.490 1.150 ;
        RECT 567.430 0.770 567.810 1.150 ;
        RECT 569.750 0.770 570.130 1.150 ;
        RECT 570.750 0.770 571.130 1.150 ;
        RECT 571.410 0.770 571.790 1.150 ;
        RECT 572.070 0.770 572.450 1.150 ;
        RECT 572.990 0.770 573.370 1.150 ;
        RECT 573.650 0.770 574.030 1.150 ;
        RECT 574.310 0.770 574.690 1.150 ;
        RECT 575.230 0.770 575.610 1.150 ;
        RECT 575.890 0.770 576.270 1.150 ;
        RECT 576.550 0.770 576.930 1.150 ;
        RECT 577.470 0.770 577.850 1.150 ;
        RECT 578.130 0.770 578.510 1.150 ;
        RECT 578.790 0.770 579.170 1.150 ;
        RECT 579.710 0.770 580.090 1.150 ;
        RECT 580.370 0.770 580.750 1.150 ;
        RECT 581.030 0.770 581.410 1.150 ;
        RECT 581.950 0.770 582.330 1.150 ;
        RECT 582.610 0.770 582.990 1.150 ;
        RECT 583.270 0.770 583.650 1.150 ;
        RECT 584.190 0.770 584.570 1.150 ;
        RECT 584.850 0.770 585.230 1.150 ;
        RECT 585.510 0.770 585.890 1.150 ;
        RECT 586.430 0.770 586.810 1.150 ;
        RECT 587.090 0.770 587.470 1.150 ;
        RECT 587.750 0.770 588.130 1.150 ;
        RECT 588.670 0.770 589.050 1.150 ;
        RECT 589.330 0.770 589.710 1.150 ;
        RECT 589.990 0.770 590.370 1.150 ;
        RECT 591.030 0.770 591.410 1.150 ;
        RECT 592.030 0.770 592.410 1.150 ;
        RECT 592.690 0.770 593.070 1.150 ;
        RECT 593.350 0.770 593.730 1.150 ;
        RECT 594.270 0.770 594.650 1.150 ;
        RECT 594.930 0.770 595.310 1.150 ;
        RECT 595.590 0.770 595.970 1.150 ;
        RECT 596.510 0.770 596.890 1.150 ;
        RECT 597.170 0.770 597.550 1.150 ;
        RECT 597.830 0.770 598.210 1.150 ;
        RECT 598.750 0.770 599.130 1.150 ;
        RECT 599.410 0.770 599.790 1.150 ;
        RECT 600.070 0.770 600.450 1.150 ;
        RECT 600.990 0.770 601.370 1.150 ;
        RECT 601.650 0.770 602.030 1.150 ;
        RECT 602.310 0.770 602.690 1.150 ;
        RECT 603.230 0.770 603.610 1.150 ;
        RECT 603.890 0.770 604.270 1.150 ;
        RECT 604.550 0.770 604.930 1.150 ;
        RECT 605.470 0.770 605.850 1.150 ;
        RECT 606.130 0.770 606.510 1.150 ;
        RECT 606.790 0.770 607.170 1.150 ;
        RECT 607.550 0.770 607.930 1.150 ;
        RECT 608.870 0.770 609.250 1.150 ;
        RECT 611.190 0.770 611.570 1.150 ;
        RECT 612.190 0.770 612.570 1.150 ;
        RECT 612.850 0.770 613.230 1.150 ;
        RECT 613.510 0.770 613.890 1.150 ;
        RECT 614.430 0.770 614.810 1.150 ;
        RECT 615.090 0.770 615.470 1.150 ;
        RECT 615.750 0.770 616.130 1.150 ;
        RECT 616.670 0.770 617.050 1.150 ;
        RECT 617.330 0.770 617.710 1.150 ;
        RECT 617.990 0.770 618.370 1.150 ;
        RECT 618.910 0.770 619.290 1.150 ;
        RECT 619.570 0.770 619.950 1.150 ;
        RECT 620.230 0.770 620.610 1.150 ;
        RECT 621.150 0.770 621.530 1.150 ;
        RECT 621.810 0.770 622.190 1.150 ;
        RECT 622.470 0.770 622.850 1.150 ;
        RECT 623.390 0.770 623.770 1.150 ;
        RECT 624.050 0.770 624.430 1.150 ;
        RECT 624.710 0.770 625.090 1.150 ;
        RECT 625.630 0.770 626.010 1.150 ;
        RECT 626.290 0.770 626.670 1.150 ;
        RECT 626.950 0.770 627.330 1.150 ;
        RECT 627.870 0.770 628.250 1.150 ;
        RECT 628.530 0.770 628.910 1.150 ;
        RECT 629.190 0.770 629.570 1.150 ;
        RECT 630.110 0.770 630.490 1.150 ;
        RECT 630.770 0.770 631.150 1.150 ;
        RECT 631.430 0.770 631.810 1.150 ;
        RECT 632.470 0.770 632.850 1.150 ;
        RECT 633.470 0.770 633.850 1.150 ;
        RECT 634.130 0.770 634.510 1.150 ;
        RECT 634.790 0.770 635.170 1.150 ;
        RECT 635.710 0.770 636.090 1.150 ;
        RECT 636.370 0.770 636.750 1.150 ;
        RECT 637.030 0.770 637.410 1.150 ;
        RECT 637.950 0.770 638.330 1.150 ;
        RECT 638.610 0.770 638.990 1.150 ;
        RECT 639.270 0.770 639.650 1.150 ;
        RECT 640.190 0.770 640.570 1.150 ;
        RECT 640.850 0.770 641.230 1.150 ;
        RECT 641.510 0.770 641.890 1.150 ;
        RECT 642.430 0.770 642.810 1.150 ;
        RECT 643.090 0.770 643.470 1.150 ;
        RECT 643.750 0.770 644.130 1.150 ;
        RECT 644.670 0.770 645.050 1.150 ;
        RECT 645.330 0.770 645.710 1.150 ;
        RECT 645.990 0.770 646.370 1.150 ;
        RECT 646.910 0.770 647.290 1.150 ;
        RECT 647.570 0.770 647.950 1.150 ;
        RECT 648.230 0.770 648.610 1.150 ;
        RECT 649.150 0.770 649.530 1.150 ;
        RECT 649.810 0.770 650.190 1.150 ;
        RECT 650.470 0.770 650.850 1.150 ;
        RECT 651.230 0.770 651.610 1.150 ;
        RECT 652.550 0.770 652.930 1.150 ;
        RECT 654.870 0.770 655.250 1.150 ;
        RECT 655.870 0.770 656.250 1.150 ;
        RECT 656.530 0.770 656.910 1.150 ;
        RECT 657.190 0.770 657.570 1.150 ;
        RECT 658.110 0.770 658.490 1.150 ;
        RECT 658.770 0.770 659.150 1.150 ;
        RECT 659.430 0.770 659.810 1.150 ;
        RECT 660.350 0.770 660.730 1.150 ;
        RECT 661.010 0.770 661.390 1.150 ;
        RECT 661.670 0.770 662.050 1.150 ;
        RECT 662.590 0.770 662.970 1.150 ;
        RECT 663.250 0.770 663.630 1.150 ;
        RECT 663.910 0.770 664.290 1.150 ;
        RECT 664.830 0.770 665.210 1.150 ;
        RECT 665.490 0.770 665.870 1.150 ;
        RECT 666.150 0.770 666.530 1.150 ;
        RECT 667.070 0.770 667.450 1.150 ;
        RECT 667.730 0.770 668.110 1.150 ;
        RECT 668.390 0.770 668.770 1.150 ;
        RECT 669.310 0.770 669.690 1.150 ;
        RECT 669.970 0.770 670.350 1.150 ;
        RECT 670.630 0.770 671.010 1.150 ;
        RECT 671.550 0.770 671.930 1.150 ;
        RECT 672.210 0.770 672.590 1.150 ;
        RECT 672.870 0.770 673.250 1.150 ;
        RECT 673.790 0.770 674.170 1.150 ;
        RECT 674.450 0.770 674.830 1.150 ;
        RECT 675.110 0.770 675.490 1.150 ;
        RECT 676.150 0.770 676.530 1.150 ;
        RECT 677.150 0.770 677.530 1.150 ;
        RECT 677.810 0.770 678.190 1.150 ;
        RECT 678.470 0.770 678.850 1.150 ;
        RECT 679.490 0.770 679.870 1.150 ;
      LAYER Via3 ;
        RECT 0.815 58.795 1.095 59.075 ;
        RECT 11.105 58.795 11.385 59.075 ;
        RECT 21.390 58.795 21.670 59.075 ;
        RECT 31.680 58.795 31.960 59.075 ;
        RECT 41.965 58.795 42.245 59.075 ;
        RECT 43.385 58.795 43.665 59.075 ;
        RECT 53.675 58.795 53.955 59.075 ;
        RECT 63.960 58.795 64.240 59.075 ;
        RECT 74.250 58.795 74.530 59.075 ;
        RECT 84.535 58.795 84.815 59.075 ;
        RECT 85.955 58.795 86.235 59.075 ;
        RECT 96.245 58.795 96.525 59.075 ;
        RECT 106.530 58.795 106.810 59.075 ;
        RECT 116.820 58.795 117.100 59.075 ;
        RECT 127.105 58.795 127.385 59.075 ;
        RECT 128.525 58.795 128.805 59.075 ;
        RECT 138.815 58.795 139.095 59.075 ;
        RECT 149.100 58.795 149.380 59.075 ;
        RECT 159.390 58.795 159.670 59.075 ;
        RECT 169.675 58.795 169.955 59.075 ;
        RECT 171.095 58.795 171.375 59.075 ;
        RECT 181.385 58.795 181.665 59.075 ;
        RECT 191.670 58.795 191.950 59.075 ;
        RECT 201.960 58.795 202.240 59.075 ;
        RECT 212.245 58.795 212.525 59.075 ;
        RECT 213.665 58.795 213.945 59.075 ;
        RECT 223.955 58.795 224.235 59.075 ;
        RECT 234.240 58.795 234.520 59.075 ;
        RECT 244.530 58.795 244.810 59.075 ;
        RECT 254.815 58.795 255.095 59.075 ;
        RECT 256.235 58.795 256.515 59.075 ;
        RECT 266.525 58.795 266.805 59.075 ;
        RECT 276.810 58.795 277.090 59.075 ;
        RECT 287.100 58.795 287.380 59.075 ;
        RECT 297.385 58.795 297.665 59.075 ;
        RECT 298.805 58.795 299.085 59.075 ;
        RECT 309.095 58.795 309.375 59.075 ;
        RECT 319.380 58.795 319.660 59.075 ;
        RECT 329.670 58.795 329.950 59.075 ;
        RECT 339.955 58.795 340.235 59.075 ;
        RECT 341.375 58.795 341.655 59.075 ;
        RECT 351.665 58.795 351.945 59.075 ;
        RECT 361.950 58.795 362.230 59.075 ;
        RECT 372.240 58.795 372.520 59.075 ;
        RECT 382.525 58.795 382.805 59.075 ;
        RECT 383.945 58.795 384.225 59.075 ;
        RECT 394.235 58.795 394.515 59.075 ;
        RECT 404.520 58.795 404.800 59.075 ;
        RECT 414.810 58.795 415.090 59.075 ;
        RECT 425.095 58.795 425.375 59.075 ;
        RECT 426.515 58.795 426.795 59.075 ;
        RECT 436.805 58.795 437.085 59.075 ;
        RECT 447.090 58.795 447.370 59.075 ;
        RECT 457.380 58.795 457.660 59.075 ;
        RECT 467.665 58.795 467.945 59.075 ;
        RECT 469.085 58.795 469.365 59.075 ;
        RECT 479.375 58.795 479.655 59.075 ;
        RECT 489.660 58.795 489.940 59.075 ;
        RECT 499.950 58.795 500.230 59.075 ;
        RECT 510.235 58.795 510.515 59.075 ;
        RECT 511.655 58.795 511.935 59.075 ;
        RECT 521.945 58.795 522.225 59.075 ;
        RECT 532.230 58.795 532.510 59.075 ;
        RECT 542.520 58.795 542.800 59.075 ;
        RECT 552.805 58.795 553.085 59.075 ;
        RECT 554.225 58.795 554.505 59.075 ;
        RECT 564.515 58.795 564.795 59.075 ;
        RECT 574.800 58.795 575.080 59.075 ;
        RECT 585.090 58.795 585.370 59.075 ;
        RECT 595.375 58.795 595.655 59.075 ;
        RECT 596.795 58.795 597.075 59.075 ;
        RECT 607.085 58.795 607.365 59.075 ;
        RECT 617.370 58.795 617.650 59.075 ;
        RECT 627.660 58.795 627.940 59.075 ;
        RECT 637.945 58.795 638.225 59.075 ;
        RECT 639.365 58.795 639.645 59.075 ;
        RECT 649.655 58.795 649.935 59.075 ;
        RECT 659.940 58.795 660.220 59.075 ;
        RECT 670.230 58.795 670.510 59.075 ;
        RECT 680.515 58.795 680.795 59.075 ;
        RECT 0.815 58.135 1.095 58.415 ;
        RECT 11.105 58.135 11.385 58.415 ;
        RECT 21.390 58.135 21.670 58.415 ;
        RECT 31.680 58.135 31.960 58.415 ;
        RECT 41.965 58.135 42.245 58.415 ;
        RECT 43.385 58.135 43.665 58.415 ;
        RECT 53.675 58.135 53.955 58.415 ;
        RECT 63.960 58.135 64.240 58.415 ;
        RECT 74.250 58.135 74.530 58.415 ;
        RECT 84.535 58.135 84.815 58.415 ;
        RECT 85.955 58.135 86.235 58.415 ;
        RECT 96.245 58.135 96.525 58.415 ;
        RECT 106.530 58.135 106.810 58.415 ;
        RECT 116.820 58.135 117.100 58.415 ;
        RECT 127.105 58.135 127.385 58.415 ;
        RECT 128.525 58.135 128.805 58.415 ;
        RECT 138.815 58.135 139.095 58.415 ;
        RECT 149.100 58.135 149.380 58.415 ;
        RECT 159.390 58.135 159.670 58.415 ;
        RECT 169.675 58.135 169.955 58.415 ;
        RECT 171.095 58.135 171.375 58.415 ;
        RECT 181.385 58.135 181.665 58.415 ;
        RECT 191.670 58.135 191.950 58.415 ;
        RECT 201.960 58.135 202.240 58.415 ;
        RECT 212.245 58.135 212.525 58.415 ;
        RECT 213.665 58.135 213.945 58.415 ;
        RECT 223.955 58.135 224.235 58.415 ;
        RECT 234.240 58.135 234.520 58.415 ;
        RECT 244.530 58.135 244.810 58.415 ;
        RECT 254.815 58.135 255.095 58.415 ;
        RECT 256.235 58.135 256.515 58.415 ;
        RECT 266.525 58.135 266.805 58.415 ;
        RECT 276.810 58.135 277.090 58.415 ;
        RECT 287.100 58.135 287.380 58.415 ;
        RECT 297.385 58.135 297.665 58.415 ;
        RECT 298.805 58.135 299.085 58.415 ;
        RECT 309.095 58.135 309.375 58.415 ;
        RECT 319.380 58.135 319.660 58.415 ;
        RECT 329.670 58.135 329.950 58.415 ;
        RECT 339.955 58.135 340.235 58.415 ;
        RECT 341.375 58.135 341.655 58.415 ;
        RECT 351.665 58.135 351.945 58.415 ;
        RECT 361.950 58.135 362.230 58.415 ;
        RECT 372.240 58.135 372.520 58.415 ;
        RECT 382.525 58.135 382.805 58.415 ;
        RECT 383.945 58.135 384.225 58.415 ;
        RECT 394.235 58.135 394.515 58.415 ;
        RECT 404.520 58.135 404.800 58.415 ;
        RECT 414.810 58.135 415.090 58.415 ;
        RECT 425.095 58.135 425.375 58.415 ;
        RECT 426.515 58.135 426.795 58.415 ;
        RECT 436.805 58.135 437.085 58.415 ;
        RECT 447.090 58.135 447.370 58.415 ;
        RECT 457.380 58.135 457.660 58.415 ;
        RECT 467.665 58.135 467.945 58.415 ;
        RECT 469.085 58.135 469.365 58.415 ;
        RECT 479.375 58.135 479.655 58.415 ;
        RECT 489.660 58.135 489.940 58.415 ;
        RECT 499.950 58.135 500.230 58.415 ;
        RECT 510.235 58.135 510.515 58.415 ;
        RECT 511.655 58.135 511.935 58.415 ;
        RECT 521.945 58.135 522.225 58.415 ;
        RECT 532.230 58.135 532.510 58.415 ;
        RECT 542.520 58.135 542.800 58.415 ;
        RECT 552.805 58.135 553.085 58.415 ;
        RECT 554.225 58.135 554.505 58.415 ;
        RECT 564.515 58.135 564.795 58.415 ;
        RECT 574.800 58.135 575.080 58.415 ;
        RECT 585.090 58.135 585.370 58.415 ;
        RECT 595.375 58.135 595.655 58.415 ;
        RECT 596.795 58.135 597.075 58.415 ;
        RECT 607.085 58.135 607.365 58.415 ;
        RECT 617.370 58.135 617.650 58.415 ;
        RECT 627.660 58.135 627.940 58.415 ;
        RECT 637.945 58.135 638.225 58.415 ;
        RECT 639.365 58.135 639.645 58.415 ;
        RECT 649.655 58.135 649.935 58.415 ;
        RECT 659.940 58.135 660.220 58.415 ;
        RECT 670.230 58.135 670.510 58.415 ;
        RECT 680.515 58.135 680.795 58.415 ;
        RECT 0.815 57.475 1.095 57.755 ;
        RECT 11.105 57.475 11.385 57.755 ;
        RECT 21.390 57.475 21.670 57.755 ;
        RECT 31.680 57.475 31.960 57.755 ;
        RECT 41.965 57.475 42.245 57.755 ;
        RECT 43.385 57.475 43.665 57.755 ;
        RECT 53.675 57.475 53.955 57.755 ;
        RECT 63.960 57.475 64.240 57.755 ;
        RECT 74.250 57.475 74.530 57.755 ;
        RECT 84.535 57.475 84.815 57.755 ;
        RECT 85.955 57.475 86.235 57.755 ;
        RECT 96.245 57.475 96.525 57.755 ;
        RECT 106.530 57.475 106.810 57.755 ;
        RECT 116.820 57.475 117.100 57.755 ;
        RECT 127.105 57.475 127.385 57.755 ;
        RECT 128.525 57.475 128.805 57.755 ;
        RECT 138.815 57.475 139.095 57.755 ;
        RECT 149.100 57.475 149.380 57.755 ;
        RECT 159.390 57.475 159.670 57.755 ;
        RECT 169.675 57.475 169.955 57.755 ;
        RECT 171.095 57.475 171.375 57.755 ;
        RECT 181.385 57.475 181.665 57.755 ;
        RECT 191.670 57.475 191.950 57.755 ;
        RECT 201.960 57.475 202.240 57.755 ;
        RECT 212.245 57.475 212.525 57.755 ;
        RECT 213.665 57.475 213.945 57.755 ;
        RECT 223.955 57.475 224.235 57.755 ;
        RECT 234.240 57.475 234.520 57.755 ;
        RECT 244.530 57.475 244.810 57.755 ;
        RECT 254.815 57.475 255.095 57.755 ;
        RECT 256.235 57.475 256.515 57.755 ;
        RECT 266.525 57.475 266.805 57.755 ;
        RECT 276.810 57.475 277.090 57.755 ;
        RECT 287.100 57.475 287.380 57.755 ;
        RECT 297.385 57.475 297.665 57.755 ;
        RECT 298.805 57.475 299.085 57.755 ;
        RECT 309.095 57.475 309.375 57.755 ;
        RECT 319.380 57.475 319.660 57.755 ;
        RECT 329.670 57.475 329.950 57.755 ;
        RECT 339.955 57.475 340.235 57.755 ;
        RECT 341.375 57.475 341.655 57.755 ;
        RECT 351.665 57.475 351.945 57.755 ;
        RECT 361.950 57.475 362.230 57.755 ;
        RECT 372.240 57.475 372.520 57.755 ;
        RECT 382.525 57.475 382.805 57.755 ;
        RECT 383.945 57.475 384.225 57.755 ;
        RECT 394.235 57.475 394.515 57.755 ;
        RECT 404.520 57.475 404.800 57.755 ;
        RECT 414.810 57.475 415.090 57.755 ;
        RECT 425.095 57.475 425.375 57.755 ;
        RECT 426.515 57.475 426.795 57.755 ;
        RECT 436.805 57.475 437.085 57.755 ;
        RECT 447.090 57.475 447.370 57.755 ;
        RECT 457.380 57.475 457.660 57.755 ;
        RECT 467.665 57.475 467.945 57.755 ;
        RECT 469.085 57.475 469.365 57.755 ;
        RECT 479.375 57.475 479.655 57.755 ;
        RECT 489.660 57.475 489.940 57.755 ;
        RECT 499.950 57.475 500.230 57.755 ;
        RECT 510.235 57.475 510.515 57.755 ;
        RECT 511.655 57.475 511.935 57.755 ;
        RECT 521.945 57.475 522.225 57.755 ;
        RECT 532.230 57.475 532.510 57.755 ;
        RECT 542.520 57.475 542.800 57.755 ;
        RECT 552.805 57.475 553.085 57.755 ;
        RECT 554.225 57.475 554.505 57.755 ;
        RECT 564.515 57.475 564.795 57.755 ;
        RECT 574.800 57.475 575.080 57.755 ;
        RECT 585.090 57.475 585.370 57.755 ;
        RECT 595.375 57.475 595.655 57.755 ;
        RECT 596.795 57.475 597.075 57.755 ;
        RECT 607.085 57.475 607.365 57.755 ;
        RECT 617.370 57.475 617.650 57.755 ;
        RECT 627.660 57.475 627.940 57.755 ;
        RECT 637.945 57.475 638.225 57.755 ;
        RECT 639.365 57.475 639.645 57.755 ;
        RECT 649.655 57.475 649.935 57.755 ;
        RECT 659.940 57.475 660.220 57.755 ;
        RECT 670.230 57.475 670.510 57.755 ;
        RECT 680.515 57.475 680.795 57.755 ;
        RECT 0.815 56.815 1.095 57.095 ;
        RECT 11.105 56.815 11.385 57.095 ;
        RECT 21.390 56.815 21.670 57.095 ;
        RECT 31.680 56.815 31.960 57.095 ;
        RECT 41.965 56.815 42.245 57.095 ;
        RECT 43.385 56.815 43.665 57.095 ;
        RECT 53.675 56.815 53.955 57.095 ;
        RECT 63.960 56.815 64.240 57.095 ;
        RECT 74.250 56.815 74.530 57.095 ;
        RECT 84.535 56.815 84.815 57.095 ;
        RECT 85.955 56.815 86.235 57.095 ;
        RECT 96.245 56.815 96.525 57.095 ;
        RECT 106.530 56.815 106.810 57.095 ;
        RECT 116.820 56.815 117.100 57.095 ;
        RECT 127.105 56.815 127.385 57.095 ;
        RECT 128.525 56.815 128.805 57.095 ;
        RECT 138.815 56.815 139.095 57.095 ;
        RECT 149.100 56.815 149.380 57.095 ;
        RECT 159.390 56.815 159.670 57.095 ;
        RECT 169.675 56.815 169.955 57.095 ;
        RECT 171.095 56.815 171.375 57.095 ;
        RECT 181.385 56.815 181.665 57.095 ;
        RECT 191.670 56.815 191.950 57.095 ;
        RECT 201.960 56.815 202.240 57.095 ;
        RECT 212.245 56.815 212.525 57.095 ;
        RECT 213.665 56.815 213.945 57.095 ;
        RECT 223.955 56.815 224.235 57.095 ;
        RECT 234.240 56.815 234.520 57.095 ;
        RECT 244.530 56.815 244.810 57.095 ;
        RECT 254.815 56.815 255.095 57.095 ;
        RECT 256.235 56.815 256.515 57.095 ;
        RECT 266.525 56.815 266.805 57.095 ;
        RECT 276.810 56.815 277.090 57.095 ;
        RECT 287.100 56.815 287.380 57.095 ;
        RECT 297.385 56.815 297.665 57.095 ;
        RECT 298.805 56.815 299.085 57.095 ;
        RECT 309.095 56.815 309.375 57.095 ;
        RECT 319.380 56.815 319.660 57.095 ;
        RECT 329.670 56.815 329.950 57.095 ;
        RECT 339.955 56.815 340.235 57.095 ;
        RECT 341.375 56.815 341.655 57.095 ;
        RECT 351.665 56.815 351.945 57.095 ;
        RECT 361.950 56.815 362.230 57.095 ;
        RECT 372.240 56.815 372.520 57.095 ;
        RECT 382.525 56.815 382.805 57.095 ;
        RECT 383.945 56.815 384.225 57.095 ;
        RECT 394.235 56.815 394.515 57.095 ;
        RECT 404.520 56.815 404.800 57.095 ;
        RECT 414.810 56.815 415.090 57.095 ;
        RECT 425.095 56.815 425.375 57.095 ;
        RECT 426.515 56.815 426.795 57.095 ;
        RECT 436.805 56.815 437.085 57.095 ;
        RECT 447.090 56.815 447.370 57.095 ;
        RECT 457.380 56.815 457.660 57.095 ;
        RECT 467.665 56.815 467.945 57.095 ;
        RECT 469.085 56.815 469.365 57.095 ;
        RECT 479.375 56.815 479.655 57.095 ;
        RECT 489.660 56.815 489.940 57.095 ;
        RECT 499.950 56.815 500.230 57.095 ;
        RECT 510.235 56.815 510.515 57.095 ;
        RECT 511.655 56.815 511.935 57.095 ;
        RECT 521.945 56.815 522.225 57.095 ;
        RECT 532.230 56.815 532.510 57.095 ;
        RECT 542.520 56.815 542.800 57.095 ;
        RECT 552.805 56.815 553.085 57.095 ;
        RECT 554.225 56.815 554.505 57.095 ;
        RECT 564.515 56.815 564.795 57.095 ;
        RECT 574.800 56.815 575.080 57.095 ;
        RECT 585.090 56.815 585.370 57.095 ;
        RECT 595.375 56.815 595.655 57.095 ;
        RECT 596.795 56.815 597.075 57.095 ;
        RECT 607.085 56.815 607.365 57.095 ;
        RECT 617.370 56.815 617.650 57.095 ;
        RECT 627.660 56.815 627.940 57.095 ;
        RECT 637.945 56.815 638.225 57.095 ;
        RECT 639.365 56.815 639.645 57.095 ;
        RECT 649.655 56.815 649.935 57.095 ;
        RECT 659.940 56.815 660.220 57.095 ;
        RECT 670.230 56.815 670.510 57.095 ;
        RECT 680.515 56.815 680.795 57.095 ;
        RECT 0.815 56.155 1.095 56.435 ;
        RECT 11.105 56.155 11.385 56.435 ;
        RECT 21.390 56.155 21.670 56.435 ;
        RECT 31.680 56.155 31.960 56.435 ;
        RECT 41.965 56.155 42.245 56.435 ;
        RECT 43.385 56.155 43.665 56.435 ;
        RECT 53.675 56.155 53.955 56.435 ;
        RECT 63.960 56.155 64.240 56.435 ;
        RECT 74.250 56.155 74.530 56.435 ;
        RECT 84.535 56.155 84.815 56.435 ;
        RECT 85.955 56.155 86.235 56.435 ;
        RECT 96.245 56.155 96.525 56.435 ;
        RECT 106.530 56.155 106.810 56.435 ;
        RECT 116.820 56.155 117.100 56.435 ;
        RECT 127.105 56.155 127.385 56.435 ;
        RECT 128.525 56.155 128.805 56.435 ;
        RECT 138.815 56.155 139.095 56.435 ;
        RECT 149.100 56.155 149.380 56.435 ;
        RECT 159.390 56.155 159.670 56.435 ;
        RECT 169.675 56.155 169.955 56.435 ;
        RECT 171.095 56.155 171.375 56.435 ;
        RECT 181.385 56.155 181.665 56.435 ;
        RECT 191.670 56.155 191.950 56.435 ;
        RECT 201.960 56.155 202.240 56.435 ;
        RECT 212.245 56.155 212.525 56.435 ;
        RECT 213.665 56.155 213.945 56.435 ;
        RECT 223.955 56.155 224.235 56.435 ;
        RECT 234.240 56.155 234.520 56.435 ;
        RECT 244.530 56.155 244.810 56.435 ;
        RECT 254.815 56.155 255.095 56.435 ;
        RECT 256.235 56.155 256.515 56.435 ;
        RECT 266.525 56.155 266.805 56.435 ;
        RECT 276.810 56.155 277.090 56.435 ;
        RECT 287.100 56.155 287.380 56.435 ;
        RECT 297.385 56.155 297.665 56.435 ;
        RECT 298.805 56.155 299.085 56.435 ;
        RECT 309.095 56.155 309.375 56.435 ;
        RECT 319.380 56.155 319.660 56.435 ;
        RECT 329.670 56.155 329.950 56.435 ;
        RECT 339.955 56.155 340.235 56.435 ;
        RECT 341.375 56.155 341.655 56.435 ;
        RECT 351.665 56.155 351.945 56.435 ;
        RECT 361.950 56.155 362.230 56.435 ;
        RECT 372.240 56.155 372.520 56.435 ;
        RECT 382.525 56.155 382.805 56.435 ;
        RECT 383.945 56.155 384.225 56.435 ;
        RECT 394.235 56.155 394.515 56.435 ;
        RECT 404.520 56.155 404.800 56.435 ;
        RECT 414.810 56.155 415.090 56.435 ;
        RECT 425.095 56.155 425.375 56.435 ;
        RECT 426.515 56.155 426.795 56.435 ;
        RECT 436.805 56.155 437.085 56.435 ;
        RECT 447.090 56.155 447.370 56.435 ;
        RECT 457.380 56.155 457.660 56.435 ;
        RECT 467.665 56.155 467.945 56.435 ;
        RECT 469.085 56.155 469.365 56.435 ;
        RECT 479.375 56.155 479.655 56.435 ;
        RECT 489.660 56.155 489.940 56.435 ;
        RECT 499.950 56.155 500.230 56.435 ;
        RECT 510.235 56.155 510.515 56.435 ;
        RECT 511.655 56.155 511.935 56.435 ;
        RECT 521.945 56.155 522.225 56.435 ;
        RECT 532.230 56.155 532.510 56.435 ;
        RECT 542.520 56.155 542.800 56.435 ;
        RECT 552.805 56.155 553.085 56.435 ;
        RECT 554.225 56.155 554.505 56.435 ;
        RECT 564.515 56.155 564.795 56.435 ;
        RECT 574.800 56.155 575.080 56.435 ;
        RECT 585.090 56.155 585.370 56.435 ;
        RECT 595.375 56.155 595.655 56.435 ;
        RECT 596.795 56.155 597.075 56.435 ;
        RECT 607.085 56.155 607.365 56.435 ;
        RECT 617.370 56.155 617.650 56.435 ;
        RECT 627.660 56.155 627.940 56.435 ;
        RECT 637.945 56.155 638.225 56.435 ;
        RECT 639.365 56.155 639.645 56.435 ;
        RECT 649.655 56.155 649.935 56.435 ;
        RECT 659.940 56.155 660.220 56.435 ;
        RECT 670.230 56.155 670.510 56.435 ;
        RECT 680.515 56.155 680.795 56.435 ;
        RECT 0.815 55.495 1.095 55.775 ;
        RECT 11.105 55.495 11.385 55.775 ;
        RECT 21.390 55.495 21.670 55.775 ;
        RECT 31.680 55.495 31.960 55.775 ;
        RECT 41.965 55.495 42.245 55.775 ;
        RECT 43.385 55.495 43.665 55.775 ;
        RECT 53.675 55.495 53.955 55.775 ;
        RECT 63.960 55.495 64.240 55.775 ;
        RECT 74.250 55.495 74.530 55.775 ;
        RECT 84.535 55.495 84.815 55.775 ;
        RECT 85.955 55.495 86.235 55.775 ;
        RECT 96.245 55.495 96.525 55.775 ;
        RECT 106.530 55.495 106.810 55.775 ;
        RECT 116.820 55.495 117.100 55.775 ;
        RECT 127.105 55.495 127.385 55.775 ;
        RECT 128.525 55.495 128.805 55.775 ;
        RECT 138.815 55.495 139.095 55.775 ;
        RECT 149.100 55.495 149.380 55.775 ;
        RECT 159.390 55.495 159.670 55.775 ;
        RECT 169.675 55.495 169.955 55.775 ;
        RECT 171.095 55.495 171.375 55.775 ;
        RECT 181.385 55.495 181.665 55.775 ;
        RECT 191.670 55.495 191.950 55.775 ;
        RECT 201.960 55.495 202.240 55.775 ;
        RECT 212.245 55.495 212.525 55.775 ;
        RECT 213.665 55.495 213.945 55.775 ;
        RECT 223.955 55.495 224.235 55.775 ;
        RECT 234.240 55.495 234.520 55.775 ;
        RECT 244.530 55.495 244.810 55.775 ;
        RECT 254.815 55.495 255.095 55.775 ;
        RECT 256.235 55.495 256.515 55.775 ;
        RECT 266.525 55.495 266.805 55.775 ;
        RECT 276.810 55.495 277.090 55.775 ;
        RECT 287.100 55.495 287.380 55.775 ;
        RECT 297.385 55.495 297.665 55.775 ;
        RECT 298.805 55.495 299.085 55.775 ;
        RECT 309.095 55.495 309.375 55.775 ;
        RECT 319.380 55.495 319.660 55.775 ;
        RECT 329.670 55.495 329.950 55.775 ;
        RECT 339.955 55.495 340.235 55.775 ;
        RECT 341.375 55.495 341.655 55.775 ;
        RECT 351.665 55.495 351.945 55.775 ;
        RECT 361.950 55.495 362.230 55.775 ;
        RECT 372.240 55.495 372.520 55.775 ;
        RECT 382.525 55.495 382.805 55.775 ;
        RECT 383.945 55.495 384.225 55.775 ;
        RECT 394.235 55.495 394.515 55.775 ;
        RECT 404.520 55.495 404.800 55.775 ;
        RECT 414.810 55.495 415.090 55.775 ;
        RECT 425.095 55.495 425.375 55.775 ;
        RECT 426.515 55.495 426.795 55.775 ;
        RECT 436.805 55.495 437.085 55.775 ;
        RECT 447.090 55.495 447.370 55.775 ;
        RECT 457.380 55.495 457.660 55.775 ;
        RECT 467.665 55.495 467.945 55.775 ;
        RECT 469.085 55.495 469.365 55.775 ;
        RECT 479.375 55.495 479.655 55.775 ;
        RECT 489.660 55.495 489.940 55.775 ;
        RECT 499.950 55.495 500.230 55.775 ;
        RECT 510.235 55.495 510.515 55.775 ;
        RECT 511.655 55.495 511.935 55.775 ;
        RECT 521.945 55.495 522.225 55.775 ;
        RECT 532.230 55.495 532.510 55.775 ;
        RECT 542.520 55.495 542.800 55.775 ;
        RECT 552.805 55.495 553.085 55.775 ;
        RECT 554.225 55.495 554.505 55.775 ;
        RECT 564.515 55.495 564.795 55.775 ;
        RECT 574.800 55.495 575.080 55.775 ;
        RECT 585.090 55.495 585.370 55.775 ;
        RECT 595.375 55.495 595.655 55.775 ;
        RECT 596.795 55.495 597.075 55.775 ;
        RECT 607.085 55.495 607.365 55.775 ;
        RECT 617.370 55.495 617.650 55.775 ;
        RECT 627.660 55.495 627.940 55.775 ;
        RECT 637.945 55.495 638.225 55.775 ;
        RECT 639.365 55.495 639.645 55.775 ;
        RECT 649.655 55.495 649.935 55.775 ;
        RECT 659.940 55.495 660.220 55.775 ;
        RECT 670.230 55.495 670.510 55.775 ;
        RECT 680.515 55.495 680.795 55.775 ;
        RECT 682.360 55.165 682.640 55.445 ;
        RECT 0.815 54.835 1.095 55.115 ;
        RECT 11.105 54.835 11.385 55.115 ;
        RECT 21.390 54.835 21.670 55.115 ;
        RECT 31.680 54.835 31.960 55.115 ;
        RECT 41.965 54.835 42.245 55.115 ;
        RECT 43.385 54.835 43.665 55.115 ;
        RECT 53.675 54.835 53.955 55.115 ;
        RECT 63.960 54.835 64.240 55.115 ;
        RECT 74.250 54.835 74.530 55.115 ;
        RECT 84.535 54.835 84.815 55.115 ;
        RECT 85.955 54.835 86.235 55.115 ;
        RECT 96.245 54.835 96.525 55.115 ;
        RECT 106.530 54.835 106.810 55.115 ;
        RECT 116.820 54.835 117.100 55.115 ;
        RECT 127.105 54.835 127.385 55.115 ;
        RECT 128.525 54.835 128.805 55.115 ;
        RECT 138.815 54.835 139.095 55.115 ;
        RECT 149.100 54.835 149.380 55.115 ;
        RECT 159.390 54.835 159.670 55.115 ;
        RECT 169.675 54.835 169.955 55.115 ;
        RECT 171.095 54.835 171.375 55.115 ;
        RECT 181.385 54.835 181.665 55.115 ;
        RECT 191.670 54.835 191.950 55.115 ;
        RECT 201.960 54.835 202.240 55.115 ;
        RECT 212.245 54.835 212.525 55.115 ;
        RECT 213.665 54.835 213.945 55.115 ;
        RECT 223.955 54.835 224.235 55.115 ;
        RECT 234.240 54.835 234.520 55.115 ;
        RECT 244.530 54.835 244.810 55.115 ;
        RECT 254.815 54.835 255.095 55.115 ;
        RECT 256.235 54.835 256.515 55.115 ;
        RECT 266.525 54.835 266.805 55.115 ;
        RECT 276.810 54.835 277.090 55.115 ;
        RECT 287.100 54.835 287.380 55.115 ;
        RECT 297.385 54.835 297.665 55.115 ;
        RECT 298.805 54.835 299.085 55.115 ;
        RECT 309.095 54.835 309.375 55.115 ;
        RECT 319.380 54.835 319.660 55.115 ;
        RECT 329.670 54.835 329.950 55.115 ;
        RECT 339.955 54.835 340.235 55.115 ;
        RECT 341.375 54.835 341.655 55.115 ;
        RECT 351.665 54.835 351.945 55.115 ;
        RECT 361.950 54.835 362.230 55.115 ;
        RECT 372.240 54.835 372.520 55.115 ;
        RECT 382.525 54.835 382.805 55.115 ;
        RECT 383.945 54.835 384.225 55.115 ;
        RECT 394.235 54.835 394.515 55.115 ;
        RECT 404.520 54.835 404.800 55.115 ;
        RECT 414.810 54.835 415.090 55.115 ;
        RECT 425.095 54.835 425.375 55.115 ;
        RECT 426.515 54.835 426.795 55.115 ;
        RECT 436.805 54.835 437.085 55.115 ;
        RECT 447.090 54.835 447.370 55.115 ;
        RECT 457.380 54.835 457.660 55.115 ;
        RECT 467.665 54.835 467.945 55.115 ;
        RECT 469.085 54.835 469.365 55.115 ;
        RECT 479.375 54.835 479.655 55.115 ;
        RECT 489.660 54.835 489.940 55.115 ;
        RECT 499.950 54.835 500.230 55.115 ;
        RECT 510.235 54.835 510.515 55.115 ;
        RECT 511.655 54.835 511.935 55.115 ;
        RECT 521.945 54.835 522.225 55.115 ;
        RECT 532.230 54.835 532.510 55.115 ;
        RECT 542.520 54.835 542.800 55.115 ;
        RECT 552.805 54.835 553.085 55.115 ;
        RECT 554.225 54.835 554.505 55.115 ;
        RECT 564.515 54.835 564.795 55.115 ;
        RECT 574.800 54.835 575.080 55.115 ;
        RECT 585.090 54.835 585.370 55.115 ;
        RECT 595.375 54.835 595.655 55.115 ;
        RECT 596.795 54.835 597.075 55.115 ;
        RECT 607.085 54.835 607.365 55.115 ;
        RECT 617.370 54.835 617.650 55.115 ;
        RECT 627.660 54.835 627.940 55.115 ;
        RECT 637.945 54.835 638.225 55.115 ;
        RECT 639.365 54.835 639.645 55.115 ;
        RECT 649.655 54.835 649.935 55.115 ;
        RECT 659.940 54.835 660.220 55.115 ;
        RECT 670.230 54.835 670.510 55.115 ;
        RECT 684.145 55.165 684.425 55.445 ;
        RECT 687.000 55.165 687.280 55.445 ;
        RECT 688.785 55.165 689.065 55.445 ;
        RECT 691.640 55.165 691.920 55.445 ;
        RECT 693.425 55.165 693.705 55.445 ;
        RECT 696.280 55.165 696.560 55.445 ;
        RECT 698.065 55.165 698.345 55.445 ;
        RECT 700.920 55.165 701.200 55.445 ;
        RECT 702.705 55.165 702.985 55.445 ;
        RECT 705.560 55.165 705.840 55.445 ;
        RECT 707.345 55.165 707.625 55.445 ;
        RECT 710.200 55.165 710.480 55.445 ;
        RECT 711.985 55.165 712.265 55.445 ;
        RECT 714.840 55.165 715.120 55.445 ;
        RECT 716.625 55.165 716.905 55.445 ;
        RECT 680.515 54.835 680.795 55.115 ;
        RECT 682.360 54.505 682.640 54.785 ;
        RECT 0.815 54.175 1.095 54.455 ;
        RECT 11.105 54.175 11.385 54.455 ;
        RECT 21.390 54.175 21.670 54.455 ;
        RECT 31.680 54.175 31.960 54.455 ;
        RECT 41.965 54.175 42.245 54.455 ;
        RECT 43.385 54.175 43.665 54.455 ;
        RECT 53.675 54.175 53.955 54.455 ;
        RECT 63.960 54.175 64.240 54.455 ;
        RECT 74.250 54.175 74.530 54.455 ;
        RECT 84.535 54.175 84.815 54.455 ;
        RECT 85.955 54.175 86.235 54.455 ;
        RECT 96.245 54.175 96.525 54.455 ;
        RECT 106.530 54.175 106.810 54.455 ;
        RECT 116.820 54.175 117.100 54.455 ;
        RECT 127.105 54.175 127.385 54.455 ;
        RECT 128.525 54.175 128.805 54.455 ;
        RECT 138.815 54.175 139.095 54.455 ;
        RECT 149.100 54.175 149.380 54.455 ;
        RECT 159.390 54.175 159.670 54.455 ;
        RECT 169.675 54.175 169.955 54.455 ;
        RECT 171.095 54.175 171.375 54.455 ;
        RECT 181.385 54.175 181.665 54.455 ;
        RECT 191.670 54.175 191.950 54.455 ;
        RECT 201.960 54.175 202.240 54.455 ;
        RECT 212.245 54.175 212.525 54.455 ;
        RECT 213.665 54.175 213.945 54.455 ;
        RECT 223.955 54.175 224.235 54.455 ;
        RECT 234.240 54.175 234.520 54.455 ;
        RECT 244.530 54.175 244.810 54.455 ;
        RECT 254.815 54.175 255.095 54.455 ;
        RECT 256.235 54.175 256.515 54.455 ;
        RECT 266.525 54.175 266.805 54.455 ;
        RECT 276.810 54.175 277.090 54.455 ;
        RECT 287.100 54.175 287.380 54.455 ;
        RECT 297.385 54.175 297.665 54.455 ;
        RECT 298.805 54.175 299.085 54.455 ;
        RECT 309.095 54.175 309.375 54.455 ;
        RECT 319.380 54.175 319.660 54.455 ;
        RECT 329.670 54.175 329.950 54.455 ;
        RECT 339.955 54.175 340.235 54.455 ;
        RECT 341.375 54.175 341.655 54.455 ;
        RECT 351.665 54.175 351.945 54.455 ;
        RECT 361.950 54.175 362.230 54.455 ;
        RECT 372.240 54.175 372.520 54.455 ;
        RECT 382.525 54.175 382.805 54.455 ;
        RECT 383.945 54.175 384.225 54.455 ;
        RECT 394.235 54.175 394.515 54.455 ;
        RECT 404.520 54.175 404.800 54.455 ;
        RECT 414.810 54.175 415.090 54.455 ;
        RECT 425.095 54.175 425.375 54.455 ;
        RECT 426.515 54.175 426.795 54.455 ;
        RECT 436.805 54.175 437.085 54.455 ;
        RECT 447.090 54.175 447.370 54.455 ;
        RECT 457.380 54.175 457.660 54.455 ;
        RECT 467.665 54.175 467.945 54.455 ;
        RECT 469.085 54.175 469.365 54.455 ;
        RECT 479.375 54.175 479.655 54.455 ;
        RECT 489.660 54.175 489.940 54.455 ;
        RECT 499.950 54.175 500.230 54.455 ;
        RECT 510.235 54.175 510.515 54.455 ;
        RECT 511.655 54.175 511.935 54.455 ;
        RECT 521.945 54.175 522.225 54.455 ;
        RECT 532.230 54.175 532.510 54.455 ;
        RECT 542.520 54.175 542.800 54.455 ;
        RECT 552.805 54.175 553.085 54.455 ;
        RECT 554.225 54.175 554.505 54.455 ;
        RECT 564.515 54.175 564.795 54.455 ;
        RECT 574.800 54.175 575.080 54.455 ;
        RECT 585.090 54.175 585.370 54.455 ;
        RECT 595.375 54.175 595.655 54.455 ;
        RECT 596.795 54.175 597.075 54.455 ;
        RECT 607.085 54.175 607.365 54.455 ;
        RECT 617.370 54.175 617.650 54.455 ;
        RECT 627.660 54.175 627.940 54.455 ;
        RECT 637.945 54.175 638.225 54.455 ;
        RECT 639.365 54.175 639.645 54.455 ;
        RECT 649.655 54.175 649.935 54.455 ;
        RECT 659.940 54.175 660.220 54.455 ;
        RECT 670.230 54.175 670.510 54.455 ;
        RECT 684.145 54.505 684.425 54.785 ;
        RECT 687.000 54.505 687.280 54.785 ;
        RECT 688.785 54.505 689.065 54.785 ;
        RECT 691.640 54.505 691.920 54.785 ;
        RECT 693.425 54.505 693.705 54.785 ;
        RECT 696.280 54.505 696.560 54.785 ;
        RECT 698.065 54.505 698.345 54.785 ;
        RECT 700.920 54.505 701.200 54.785 ;
        RECT 702.705 54.505 702.985 54.785 ;
        RECT 705.560 54.505 705.840 54.785 ;
        RECT 707.345 54.505 707.625 54.785 ;
        RECT 710.200 54.505 710.480 54.785 ;
        RECT 711.985 54.505 712.265 54.785 ;
        RECT 714.840 54.505 715.120 54.785 ;
        RECT 716.625 54.505 716.905 54.785 ;
        RECT 680.515 54.175 680.795 54.455 ;
        RECT 682.360 53.845 682.640 54.125 ;
        RECT 0.815 53.515 1.095 53.795 ;
        RECT 11.105 53.515 11.385 53.795 ;
        RECT 21.390 53.515 21.670 53.795 ;
        RECT 31.680 53.515 31.960 53.795 ;
        RECT 41.965 53.515 42.245 53.795 ;
        RECT 43.385 53.515 43.665 53.795 ;
        RECT 53.675 53.515 53.955 53.795 ;
        RECT 63.960 53.515 64.240 53.795 ;
        RECT 74.250 53.515 74.530 53.795 ;
        RECT 84.535 53.515 84.815 53.795 ;
        RECT 85.955 53.515 86.235 53.795 ;
        RECT 96.245 53.515 96.525 53.795 ;
        RECT 106.530 53.515 106.810 53.795 ;
        RECT 116.820 53.515 117.100 53.795 ;
        RECT 127.105 53.515 127.385 53.795 ;
        RECT 128.525 53.515 128.805 53.795 ;
        RECT 138.815 53.515 139.095 53.795 ;
        RECT 149.100 53.515 149.380 53.795 ;
        RECT 159.390 53.515 159.670 53.795 ;
        RECT 169.675 53.515 169.955 53.795 ;
        RECT 171.095 53.515 171.375 53.795 ;
        RECT 181.385 53.515 181.665 53.795 ;
        RECT 191.670 53.515 191.950 53.795 ;
        RECT 201.960 53.515 202.240 53.795 ;
        RECT 212.245 53.515 212.525 53.795 ;
        RECT 213.665 53.515 213.945 53.795 ;
        RECT 223.955 53.515 224.235 53.795 ;
        RECT 234.240 53.515 234.520 53.795 ;
        RECT 244.530 53.515 244.810 53.795 ;
        RECT 254.815 53.515 255.095 53.795 ;
        RECT 256.235 53.515 256.515 53.795 ;
        RECT 266.525 53.515 266.805 53.795 ;
        RECT 276.810 53.515 277.090 53.795 ;
        RECT 287.100 53.515 287.380 53.795 ;
        RECT 297.385 53.515 297.665 53.795 ;
        RECT 298.805 53.515 299.085 53.795 ;
        RECT 309.095 53.515 309.375 53.795 ;
        RECT 319.380 53.515 319.660 53.795 ;
        RECT 329.670 53.515 329.950 53.795 ;
        RECT 339.955 53.515 340.235 53.795 ;
        RECT 341.375 53.515 341.655 53.795 ;
        RECT 351.665 53.515 351.945 53.795 ;
        RECT 361.950 53.515 362.230 53.795 ;
        RECT 372.240 53.515 372.520 53.795 ;
        RECT 382.525 53.515 382.805 53.795 ;
        RECT 383.945 53.515 384.225 53.795 ;
        RECT 394.235 53.515 394.515 53.795 ;
        RECT 404.520 53.515 404.800 53.795 ;
        RECT 414.810 53.515 415.090 53.795 ;
        RECT 425.095 53.515 425.375 53.795 ;
        RECT 426.515 53.515 426.795 53.795 ;
        RECT 436.805 53.515 437.085 53.795 ;
        RECT 447.090 53.515 447.370 53.795 ;
        RECT 457.380 53.515 457.660 53.795 ;
        RECT 467.665 53.515 467.945 53.795 ;
        RECT 469.085 53.515 469.365 53.795 ;
        RECT 479.375 53.515 479.655 53.795 ;
        RECT 489.660 53.515 489.940 53.795 ;
        RECT 499.950 53.515 500.230 53.795 ;
        RECT 510.235 53.515 510.515 53.795 ;
        RECT 511.655 53.515 511.935 53.795 ;
        RECT 521.945 53.515 522.225 53.795 ;
        RECT 532.230 53.515 532.510 53.795 ;
        RECT 542.520 53.515 542.800 53.795 ;
        RECT 552.805 53.515 553.085 53.795 ;
        RECT 554.225 53.515 554.505 53.795 ;
        RECT 564.515 53.515 564.795 53.795 ;
        RECT 574.800 53.515 575.080 53.795 ;
        RECT 585.090 53.515 585.370 53.795 ;
        RECT 595.375 53.515 595.655 53.795 ;
        RECT 596.795 53.515 597.075 53.795 ;
        RECT 607.085 53.515 607.365 53.795 ;
        RECT 617.370 53.515 617.650 53.795 ;
        RECT 627.660 53.515 627.940 53.795 ;
        RECT 637.945 53.515 638.225 53.795 ;
        RECT 639.365 53.515 639.645 53.795 ;
        RECT 649.655 53.515 649.935 53.795 ;
        RECT 659.940 53.515 660.220 53.795 ;
        RECT 670.230 53.515 670.510 53.795 ;
        RECT 684.145 53.845 684.425 54.125 ;
        RECT 687.000 53.845 687.280 54.125 ;
        RECT 688.785 53.845 689.065 54.125 ;
        RECT 691.640 53.845 691.920 54.125 ;
        RECT 693.425 53.845 693.705 54.125 ;
        RECT 696.280 53.845 696.560 54.125 ;
        RECT 698.065 53.845 698.345 54.125 ;
        RECT 700.920 53.845 701.200 54.125 ;
        RECT 702.705 53.845 702.985 54.125 ;
        RECT 705.560 53.845 705.840 54.125 ;
        RECT 707.345 53.845 707.625 54.125 ;
        RECT 710.200 53.845 710.480 54.125 ;
        RECT 711.985 53.845 712.265 54.125 ;
        RECT 714.840 53.845 715.120 54.125 ;
        RECT 716.625 53.845 716.905 54.125 ;
        RECT 680.515 53.515 680.795 53.795 ;
        RECT 682.360 53.185 682.640 53.465 ;
        RECT 0.815 52.855 1.095 53.135 ;
        RECT 11.105 52.855 11.385 53.135 ;
        RECT 21.390 52.855 21.670 53.135 ;
        RECT 31.680 52.855 31.960 53.135 ;
        RECT 41.965 52.855 42.245 53.135 ;
        RECT 43.385 52.855 43.665 53.135 ;
        RECT 53.675 52.855 53.955 53.135 ;
        RECT 63.960 52.855 64.240 53.135 ;
        RECT 74.250 52.855 74.530 53.135 ;
        RECT 84.535 52.855 84.815 53.135 ;
        RECT 85.955 52.855 86.235 53.135 ;
        RECT 96.245 52.855 96.525 53.135 ;
        RECT 106.530 52.855 106.810 53.135 ;
        RECT 116.820 52.855 117.100 53.135 ;
        RECT 127.105 52.855 127.385 53.135 ;
        RECT 128.525 52.855 128.805 53.135 ;
        RECT 138.815 52.855 139.095 53.135 ;
        RECT 149.100 52.855 149.380 53.135 ;
        RECT 159.390 52.855 159.670 53.135 ;
        RECT 169.675 52.855 169.955 53.135 ;
        RECT 171.095 52.855 171.375 53.135 ;
        RECT 181.385 52.855 181.665 53.135 ;
        RECT 191.670 52.855 191.950 53.135 ;
        RECT 201.960 52.855 202.240 53.135 ;
        RECT 212.245 52.855 212.525 53.135 ;
        RECT 213.665 52.855 213.945 53.135 ;
        RECT 223.955 52.855 224.235 53.135 ;
        RECT 234.240 52.855 234.520 53.135 ;
        RECT 244.530 52.855 244.810 53.135 ;
        RECT 254.815 52.855 255.095 53.135 ;
        RECT 256.235 52.855 256.515 53.135 ;
        RECT 266.525 52.855 266.805 53.135 ;
        RECT 276.810 52.855 277.090 53.135 ;
        RECT 287.100 52.855 287.380 53.135 ;
        RECT 297.385 52.855 297.665 53.135 ;
        RECT 298.805 52.855 299.085 53.135 ;
        RECT 309.095 52.855 309.375 53.135 ;
        RECT 319.380 52.855 319.660 53.135 ;
        RECT 329.670 52.855 329.950 53.135 ;
        RECT 339.955 52.855 340.235 53.135 ;
        RECT 341.375 52.855 341.655 53.135 ;
        RECT 351.665 52.855 351.945 53.135 ;
        RECT 361.950 52.855 362.230 53.135 ;
        RECT 372.240 52.855 372.520 53.135 ;
        RECT 382.525 52.855 382.805 53.135 ;
        RECT 383.945 52.855 384.225 53.135 ;
        RECT 394.235 52.855 394.515 53.135 ;
        RECT 404.520 52.855 404.800 53.135 ;
        RECT 414.810 52.855 415.090 53.135 ;
        RECT 425.095 52.855 425.375 53.135 ;
        RECT 426.515 52.855 426.795 53.135 ;
        RECT 436.805 52.855 437.085 53.135 ;
        RECT 447.090 52.855 447.370 53.135 ;
        RECT 457.380 52.855 457.660 53.135 ;
        RECT 467.665 52.855 467.945 53.135 ;
        RECT 469.085 52.855 469.365 53.135 ;
        RECT 479.375 52.855 479.655 53.135 ;
        RECT 489.660 52.855 489.940 53.135 ;
        RECT 499.950 52.855 500.230 53.135 ;
        RECT 510.235 52.855 510.515 53.135 ;
        RECT 511.655 52.855 511.935 53.135 ;
        RECT 521.945 52.855 522.225 53.135 ;
        RECT 532.230 52.855 532.510 53.135 ;
        RECT 542.520 52.855 542.800 53.135 ;
        RECT 552.805 52.855 553.085 53.135 ;
        RECT 554.225 52.855 554.505 53.135 ;
        RECT 564.515 52.855 564.795 53.135 ;
        RECT 574.800 52.855 575.080 53.135 ;
        RECT 585.090 52.855 585.370 53.135 ;
        RECT 595.375 52.855 595.655 53.135 ;
        RECT 596.795 52.855 597.075 53.135 ;
        RECT 607.085 52.855 607.365 53.135 ;
        RECT 617.370 52.855 617.650 53.135 ;
        RECT 627.660 52.855 627.940 53.135 ;
        RECT 637.945 52.855 638.225 53.135 ;
        RECT 639.365 52.855 639.645 53.135 ;
        RECT 649.655 52.855 649.935 53.135 ;
        RECT 659.940 52.855 660.220 53.135 ;
        RECT 670.230 52.855 670.510 53.135 ;
        RECT 684.145 53.185 684.425 53.465 ;
        RECT 687.000 53.185 687.280 53.465 ;
        RECT 688.785 53.185 689.065 53.465 ;
        RECT 691.640 53.185 691.920 53.465 ;
        RECT 693.425 53.185 693.705 53.465 ;
        RECT 696.280 53.185 696.560 53.465 ;
        RECT 698.065 53.185 698.345 53.465 ;
        RECT 700.920 53.185 701.200 53.465 ;
        RECT 702.705 53.185 702.985 53.465 ;
        RECT 705.560 53.185 705.840 53.465 ;
        RECT 707.345 53.185 707.625 53.465 ;
        RECT 710.200 53.185 710.480 53.465 ;
        RECT 711.985 53.185 712.265 53.465 ;
        RECT 714.840 53.185 715.120 53.465 ;
        RECT 716.625 53.185 716.905 53.465 ;
        RECT 680.515 52.855 680.795 53.135 ;
        RECT 682.360 52.525 682.640 52.805 ;
        RECT 0.815 52.195 1.095 52.475 ;
        RECT 11.105 52.195 11.385 52.475 ;
        RECT 21.390 52.195 21.670 52.475 ;
        RECT 31.680 52.195 31.960 52.475 ;
        RECT 41.965 52.195 42.245 52.475 ;
        RECT 43.385 52.195 43.665 52.475 ;
        RECT 53.675 52.195 53.955 52.475 ;
        RECT 63.960 52.195 64.240 52.475 ;
        RECT 74.250 52.195 74.530 52.475 ;
        RECT 84.535 52.195 84.815 52.475 ;
        RECT 85.955 52.195 86.235 52.475 ;
        RECT 96.245 52.195 96.525 52.475 ;
        RECT 106.530 52.195 106.810 52.475 ;
        RECT 116.820 52.195 117.100 52.475 ;
        RECT 127.105 52.195 127.385 52.475 ;
        RECT 128.525 52.195 128.805 52.475 ;
        RECT 138.815 52.195 139.095 52.475 ;
        RECT 149.100 52.195 149.380 52.475 ;
        RECT 159.390 52.195 159.670 52.475 ;
        RECT 169.675 52.195 169.955 52.475 ;
        RECT 171.095 52.195 171.375 52.475 ;
        RECT 181.385 52.195 181.665 52.475 ;
        RECT 191.670 52.195 191.950 52.475 ;
        RECT 201.960 52.195 202.240 52.475 ;
        RECT 212.245 52.195 212.525 52.475 ;
        RECT 213.665 52.195 213.945 52.475 ;
        RECT 223.955 52.195 224.235 52.475 ;
        RECT 234.240 52.195 234.520 52.475 ;
        RECT 244.530 52.195 244.810 52.475 ;
        RECT 254.815 52.195 255.095 52.475 ;
        RECT 256.235 52.195 256.515 52.475 ;
        RECT 266.525 52.195 266.805 52.475 ;
        RECT 276.810 52.195 277.090 52.475 ;
        RECT 287.100 52.195 287.380 52.475 ;
        RECT 297.385 52.195 297.665 52.475 ;
        RECT 298.805 52.195 299.085 52.475 ;
        RECT 309.095 52.195 309.375 52.475 ;
        RECT 319.380 52.195 319.660 52.475 ;
        RECT 329.670 52.195 329.950 52.475 ;
        RECT 339.955 52.195 340.235 52.475 ;
        RECT 341.375 52.195 341.655 52.475 ;
        RECT 351.665 52.195 351.945 52.475 ;
        RECT 361.950 52.195 362.230 52.475 ;
        RECT 372.240 52.195 372.520 52.475 ;
        RECT 382.525 52.195 382.805 52.475 ;
        RECT 383.945 52.195 384.225 52.475 ;
        RECT 394.235 52.195 394.515 52.475 ;
        RECT 404.520 52.195 404.800 52.475 ;
        RECT 414.810 52.195 415.090 52.475 ;
        RECT 425.095 52.195 425.375 52.475 ;
        RECT 426.515 52.195 426.795 52.475 ;
        RECT 436.805 52.195 437.085 52.475 ;
        RECT 447.090 52.195 447.370 52.475 ;
        RECT 457.380 52.195 457.660 52.475 ;
        RECT 467.665 52.195 467.945 52.475 ;
        RECT 469.085 52.195 469.365 52.475 ;
        RECT 479.375 52.195 479.655 52.475 ;
        RECT 489.660 52.195 489.940 52.475 ;
        RECT 499.950 52.195 500.230 52.475 ;
        RECT 510.235 52.195 510.515 52.475 ;
        RECT 511.655 52.195 511.935 52.475 ;
        RECT 521.945 52.195 522.225 52.475 ;
        RECT 532.230 52.195 532.510 52.475 ;
        RECT 542.520 52.195 542.800 52.475 ;
        RECT 552.805 52.195 553.085 52.475 ;
        RECT 554.225 52.195 554.505 52.475 ;
        RECT 564.515 52.195 564.795 52.475 ;
        RECT 574.800 52.195 575.080 52.475 ;
        RECT 585.090 52.195 585.370 52.475 ;
        RECT 595.375 52.195 595.655 52.475 ;
        RECT 596.795 52.195 597.075 52.475 ;
        RECT 607.085 52.195 607.365 52.475 ;
        RECT 617.370 52.195 617.650 52.475 ;
        RECT 627.660 52.195 627.940 52.475 ;
        RECT 637.945 52.195 638.225 52.475 ;
        RECT 639.365 52.195 639.645 52.475 ;
        RECT 649.655 52.195 649.935 52.475 ;
        RECT 659.940 52.195 660.220 52.475 ;
        RECT 670.230 52.195 670.510 52.475 ;
        RECT 684.145 52.525 684.425 52.805 ;
        RECT 687.000 52.525 687.280 52.805 ;
        RECT 688.785 52.525 689.065 52.805 ;
        RECT 691.640 52.525 691.920 52.805 ;
        RECT 693.425 52.525 693.705 52.805 ;
        RECT 696.280 52.525 696.560 52.805 ;
        RECT 698.065 52.525 698.345 52.805 ;
        RECT 700.920 52.525 701.200 52.805 ;
        RECT 702.705 52.525 702.985 52.805 ;
        RECT 705.560 52.525 705.840 52.805 ;
        RECT 707.345 52.525 707.625 52.805 ;
        RECT 710.200 52.525 710.480 52.805 ;
        RECT 711.985 52.525 712.265 52.805 ;
        RECT 714.840 52.525 715.120 52.805 ;
        RECT 716.625 52.525 716.905 52.805 ;
        RECT 680.515 52.195 680.795 52.475 ;
        RECT 682.360 51.865 682.640 52.145 ;
        RECT 0.815 51.535 1.095 51.815 ;
        RECT 11.105 51.535 11.385 51.815 ;
        RECT 21.390 51.535 21.670 51.815 ;
        RECT 31.680 51.535 31.960 51.815 ;
        RECT 41.965 51.535 42.245 51.815 ;
        RECT 43.385 51.535 43.665 51.815 ;
        RECT 53.675 51.535 53.955 51.815 ;
        RECT 63.960 51.535 64.240 51.815 ;
        RECT 74.250 51.535 74.530 51.815 ;
        RECT 84.535 51.535 84.815 51.815 ;
        RECT 85.955 51.535 86.235 51.815 ;
        RECT 96.245 51.535 96.525 51.815 ;
        RECT 106.530 51.535 106.810 51.815 ;
        RECT 116.820 51.535 117.100 51.815 ;
        RECT 127.105 51.535 127.385 51.815 ;
        RECT 128.525 51.535 128.805 51.815 ;
        RECT 138.815 51.535 139.095 51.815 ;
        RECT 149.100 51.535 149.380 51.815 ;
        RECT 159.390 51.535 159.670 51.815 ;
        RECT 169.675 51.535 169.955 51.815 ;
        RECT 171.095 51.535 171.375 51.815 ;
        RECT 181.385 51.535 181.665 51.815 ;
        RECT 191.670 51.535 191.950 51.815 ;
        RECT 201.960 51.535 202.240 51.815 ;
        RECT 212.245 51.535 212.525 51.815 ;
        RECT 213.665 51.535 213.945 51.815 ;
        RECT 223.955 51.535 224.235 51.815 ;
        RECT 234.240 51.535 234.520 51.815 ;
        RECT 244.530 51.535 244.810 51.815 ;
        RECT 254.815 51.535 255.095 51.815 ;
        RECT 256.235 51.535 256.515 51.815 ;
        RECT 266.525 51.535 266.805 51.815 ;
        RECT 276.810 51.535 277.090 51.815 ;
        RECT 287.100 51.535 287.380 51.815 ;
        RECT 297.385 51.535 297.665 51.815 ;
        RECT 298.805 51.535 299.085 51.815 ;
        RECT 309.095 51.535 309.375 51.815 ;
        RECT 319.380 51.535 319.660 51.815 ;
        RECT 329.670 51.535 329.950 51.815 ;
        RECT 339.955 51.535 340.235 51.815 ;
        RECT 341.375 51.535 341.655 51.815 ;
        RECT 351.665 51.535 351.945 51.815 ;
        RECT 361.950 51.535 362.230 51.815 ;
        RECT 372.240 51.535 372.520 51.815 ;
        RECT 382.525 51.535 382.805 51.815 ;
        RECT 383.945 51.535 384.225 51.815 ;
        RECT 394.235 51.535 394.515 51.815 ;
        RECT 404.520 51.535 404.800 51.815 ;
        RECT 414.810 51.535 415.090 51.815 ;
        RECT 425.095 51.535 425.375 51.815 ;
        RECT 426.515 51.535 426.795 51.815 ;
        RECT 436.805 51.535 437.085 51.815 ;
        RECT 447.090 51.535 447.370 51.815 ;
        RECT 457.380 51.535 457.660 51.815 ;
        RECT 467.665 51.535 467.945 51.815 ;
        RECT 469.085 51.535 469.365 51.815 ;
        RECT 479.375 51.535 479.655 51.815 ;
        RECT 489.660 51.535 489.940 51.815 ;
        RECT 499.950 51.535 500.230 51.815 ;
        RECT 510.235 51.535 510.515 51.815 ;
        RECT 511.655 51.535 511.935 51.815 ;
        RECT 521.945 51.535 522.225 51.815 ;
        RECT 532.230 51.535 532.510 51.815 ;
        RECT 542.520 51.535 542.800 51.815 ;
        RECT 552.805 51.535 553.085 51.815 ;
        RECT 554.225 51.535 554.505 51.815 ;
        RECT 564.515 51.535 564.795 51.815 ;
        RECT 574.800 51.535 575.080 51.815 ;
        RECT 585.090 51.535 585.370 51.815 ;
        RECT 595.375 51.535 595.655 51.815 ;
        RECT 596.795 51.535 597.075 51.815 ;
        RECT 607.085 51.535 607.365 51.815 ;
        RECT 617.370 51.535 617.650 51.815 ;
        RECT 627.660 51.535 627.940 51.815 ;
        RECT 637.945 51.535 638.225 51.815 ;
        RECT 639.365 51.535 639.645 51.815 ;
        RECT 649.655 51.535 649.935 51.815 ;
        RECT 659.940 51.535 660.220 51.815 ;
        RECT 670.230 51.535 670.510 51.815 ;
        RECT 684.145 51.865 684.425 52.145 ;
        RECT 687.000 51.865 687.280 52.145 ;
        RECT 688.785 51.865 689.065 52.145 ;
        RECT 691.640 51.865 691.920 52.145 ;
        RECT 693.425 51.865 693.705 52.145 ;
        RECT 696.280 51.865 696.560 52.145 ;
        RECT 698.065 51.865 698.345 52.145 ;
        RECT 700.920 51.865 701.200 52.145 ;
        RECT 702.705 51.865 702.985 52.145 ;
        RECT 705.560 51.865 705.840 52.145 ;
        RECT 707.345 51.865 707.625 52.145 ;
        RECT 710.200 51.865 710.480 52.145 ;
        RECT 711.985 51.865 712.265 52.145 ;
        RECT 714.840 51.865 715.120 52.145 ;
        RECT 716.625 51.865 716.905 52.145 ;
        RECT 680.515 51.535 680.795 51.815 ;
        RECT 682.360 51.205 682.640 51.485 ;
        RECT 0.815 50.875 1.095 51.155 ;
        RECT 11.105 50.875 11.385 51.155 ;
        RECT 21.390 50.875 21.670 51.155 ;
        RECT 31.680 50.875 31.960 51.155 ;
        RECT 41.965 50.875 42.245 51.155 ;
        RECT 43.385 50.875 43.665 51.155 ;
        RECT 53.675 50.875 53.955 51.155 ;
        RECT 63.960 50.875 64.240 51.155 ;
        RECT 74.250 50.875 74.530 51.155 ;
        RECT 84.535 50.875 84.815 51.155 ;
        RECT 85.955 50.875 86.235 51.155 ;
        RECT 96.245 50.875 96.525 51.155 ;
        RECT 106.530 50.875 106.810 51.155 ;
        RECT 116.820 50.875 117.100 51.155 ;
        RECT 127.105 50.875 127.385 51.155 ;
        RECT 128.525 50.875 128.805 51.155 ;
        RECT 138.815 50.875 139.095 51.155 ;
        RECT 149.100 50.875 149.380 51.155 ;
        RECT 159.390 50.875 159.670 51.155 ;
        RECT 169.675 50.875 169.955 51.155 ;
        RECT 171.095 50.875 171.375 51.155 ;
        RECT 181.385 50.875 181.665 51.155 ;
        RECT 191.670 50.875 191.950 51.155 ;
        RECT 201.960 50.875 202.240 51.155 ;
        RECT 212.245 50.875 212.525 51.155 ;
        RECT 213.665 50.875 213.945 51.155 ;
        RECT 223.955 50.875 224.235 51.155 ;
        RECT 234.240 50.875 234.520 51.155 ;
        RECT 244.530 50.875 244.810 51.155 ;
        RECT 254.815 50.875 255.095 51.155 ;
        RECT 256.235 50.875 256.515 51.155 ;
        RECT 266.525 50.875 266.805 51.155 ;
        RECT 276.810 50.875 277.090 51.155 ;
        RECT 287.100 50.875 287.380 51.155 ;
        RECT 297.385 50.875 297.665 51.155 ;
        RECT 298.805 50.875 299.085 51.155 ;
        RECT 309.095 50.875 309.375 51.155 ;
        RECT 319.380 50.875 319.660 51.155 ;
        RECT 329.670 50.875 329.950 51.155 ;
        RECT 339.955 50.875 340.235 51.155 ;
        RECT 341.375 50.875 341.655 51.155 ;
        RECT 351.665 50.875 351.945 51.155 ;
        RECT 361.950 50.875 362.230 51.155 ;
        RECT 372.240 50.875 372.520 51.155 ;
        RECT 382.525 50.875 382.805 51.155 ;
        RECT 383.945 50.875 384.225 51.155 ;
        RECT 394.235 50.875 394.515 51.155 ;
        RECT 404.520 50.875 404.800 51.155 ;
        RECT 414.810 50.875 415.090 51.155 ;
        RECT 425.095 50.875 425.375 51.155 ;
        RECT 426.515 50.875 426.795 51.155 ;
        RECT 436.805 50.875 437.085 51.155 ;
        RECT 447.090 50.875 447.370 51.155 ;
        RECT 457.380 50.875 457.660 51.155 ;
        RECT 467.665 50.875 467.945 51.155 ;
        RECT 469.085 50.875 469.365 51.155 ;
        RECT 479.375 50.875 479.655 51.155 ;
        RECT 489.660 50.875 489.940 51.155 ;
        RECT 499.950 50.875 500.230 51.155 ;
        RECT 510.235 50.875 510.515 51.155 ;
        RECT 511.655 50.875 511.935 51.155 ;
        RECT 521.945 50.875 522.225 51.155 ;
        RECT 532.230 50.875 532.510 51.155 ;
        RECT 542.520 50.875 542.800 51.155 ;
        RECT 552.805 50.875 553.085 51.155 ;
        RECT 554.225 50.875 554.505 51.155 ;
        RECT 564.515 50.875 564.795 51.155 ;
        RECT 574.800 50.875 575.080 51.155 ;
        RECT 585.090 50.875 585.370 51.155 ;
        RECT 595.375 50.875 595.655 51.155 ;
        RECT 596.795 50.875 597.075 51.155 ;
        RECT 607.085 50.875 607.365 51.155 ;
        RECT 617.370 50.875 617.650 51.155 ;
        RECT 627.660 50.875 627.940 51.155 ;
        RECT 637.945 50.875 638.225 51.155 ;
        RECT 639.365 50.875 639.645 51.155 ;
        RECT 649.655 50.875 649.935 51.155 ;
        RECT 659.940 50.875 660.220 51.155 ;
        RECT 670.230 50.875 670.510 51.155 ;
        RECT 684.145 51.205 684.425 51.485 ;
        RECT 687.000 51.205 687.280 51.485 ;
        RECT 688.785 51.205 689.065 51.485 ;
        RECT 691.640 51.205 691.920 51.485 ;
        RECT 693.425 51.205 693.705 51.485 ;
        RECT 696.280 51.205 696.560 51.485 ;
        RECT 698.065 51.205 698.345 51.485 ;
        RECT 700.920 51.205 701.200 51.485 ;
        RECT 702.705 51.205 702.985 51.485 ;
        RECT 705.560 51.205 705.840 51.485 ;
        RECT 707.345 51.205 707.625 51.485 ;
        RECT 710.200 51.205 710.480 51.485 ;
        RECT 711.985 51.205 712.265 51.485 ;
        RECT 714.840 51.205 715.120 51.485 ;
        RECT 716.625 51.205 716.905 51.485 ;
        RECT 680.515 50.875 680.795 51.155 ;
        RECT 682.360 50.545 682.640 50.825 ;
        RECT 0.815 50.215 1.095 50.495 ;
        RECT 11.105 50.215 11.385 50.495 ;
        RECT 21.390 50.215 21.670 50.495 ;
        RECT 31.680 50.215 31.960 50.495 ;
        RECT 41.965 50.215 42.245 50.495 ;
        RECT 43.385 50.215 43.665 50.495 ;
        RECT 53.675 50.215 53.955 50.495 ;
        RECT 63.960 50.215 64.240 50.495 ;
        RECT 74.250 50.215 74.530 50.495 ;
        RECT 84.535 50.215 84.815 50.495 ;
        RECT 85.955 50.215 86.235 50.495 ;
        RECT 96.245 50.215 96.525 50.495 ;
        RECT 106.530 50.215 106.810 50.495 ;
        RECT 116.820 50.215 117.100 50.495 ;
        RECT 127.105 50.215 127.385 50.495 ;
        RECT 128.525 50.215 128.805 50.495 ;
        RECT 138.815 50.215 139.095 50.495 ;
        RECT 149.100 50.215 149.380 50.495 ;
        RECT 159.390 50.215 159.670 50.495 ;
        RECT 169.675 50.215 169.955 50.495 ;
        RECT 171.095 50.215 171.375 50.495 ;
        RECT 181.385 50.215 181.665 50.495 ;
        RECT 191.670 50.215 191.950 50.495 ;
        RECT 201.960 50.215 202.240 50.495 ;
        RECT 212.245 50.215 212.525 50.495 ;
        RECT 213.665 50.215 213.945 50.495 ;
        RECT 223.955 50.215 224.235 50.495 ;
        RECT 234.240 50.215 234.520 50.495 ;
        RECT 244.530 50.215 244.810 50.495 ;
        RECT 254.815 50.215 255.095 50.495 ;
        RECT 256.235 50.215 256.515 50.495 ;
        RECT 266.525 50.215 266.805 50.495 ;
        RECT 276.810 50.215 277.090 50.495 ;
        RECT 287.100 50.215 287.380 50.495 ;
        RECT 297.385 50.215 297.665 50.495 ;
        RECT 298.805 50.215 299.085 50.495 ;
        RECT 309.095 50.215 309.375 50.495 ;
        RECT 319.380 50.215 319.660 50.495 ;
        RECT 329.670 50.215 329.950 50.495 ;
        RECT 339.955 50.215 340.235 50.495 ;
        RECT 341.375 50.215 341.655 50.495 ;
        RECT 351.665 50.215 351.945 50.495 ;
        RECT 361.950 50.215 362.230 50.495 ;
        RECT 372.240 50.215 372.520 50.495 ;
        RECT 382.525 50.215 382.805 50.495 ;
        RECT 383.945 50.215 384.225 50.495 ;
        RECT 394.235 50.215 394.515 50.495 ;
        RECT 404.520 50.215 404.800 50.495 ;
        RECT 414.810 50.215 415.090 50.495 ;
        RECT 425.095 50.215 425.375 50.495 ;
        RECT 426.515 50.215 426.795 50.495 ;
        RECT 436.805 50.215 437.085 50.495 ;
        RECT 447.090 50.215 447.370 50.495 ;
        RECT 457.380 50.215 457.660 50.495 ;
        RECT 467.665 50.215 467.945 50.495 ;
        RECT 469.085 50.215 469.365 50.495 ;
        RECT 479.375 50.215 479.655 50.495 ;
        RECT 489.660 50.215 489.940 50.495 ;
        RECT 499.950 50.215 500.230 50.495 ;
        RECT 510.235 50.215 510.515 50.495 ;
        RECT 511.655 50.215 511.935 50.495 ;
        RECT 521.945 50.215 522.225 50.495 ;
        RECT 532.230 50.215 532.510 50.495 ;
        RECT 542.520 50.215 542.800 50.495 ;
        RECT 552.805 50.215 553.085 50.495 ;
        RECT 554.225 50.215 554.505 50.495 ;
        RECT 564.515 50.215 564.795 50.495 ;
        RECT 574.800 50.215 575.080 50.495 ;
        RECT 585.090 50.215 585.370 50.495 ;
        RECT 595.375 50.215 595.655 50.495 ;
        RECT 596.795 50.215 597.075 50.495 ;
        RECT 607.085 50.215 607.365 50.495 ;
        RECT 617.370 50.215 617.650 50.495 ;
        RECT 627.660 50.215 627.940 50.495 ;
        RECT 637.945 50.215 638.225 50.495 ;
        RECT 639.365 50.215 639.645 50.495 ;
        RECT 649.655 50.215 649.935 50.495 ;
        RECT 659.940 50.215 660.220 50.495 ;
        RECT 670.230 50.215 670.510 50.495 ;
        RECT 684.145 50.545 684.425 50.825 ;
        RECT 687.000 50.545 687.280 50.825 ;
        RECT 688.785 50.545 689.065 50.825 ;
        RECT 691.640 50.545 691.920 50.825 ;
        RECT 693.425 50.545 693.705 50.825 ;
        RECT 696.280 50.545 696.560 50.825 ;
        RECT 698.065 50.545 698.345 50.825 ;
        RECT 700.920 50.545 701.200 50.825 ;
        RECT 702.705 50.545 702.985 50.825 ;
        RECT 705.560 50.545 705.840 50.825 ;
        RECT 707.345 50.545 707.625 50.825 ;
        RECT 710.200 50.545 710.480 50.825 ;
        RECT 711.985 50.545 712.265 50.825 ;
        RECT 714.840 50.545 715.120 50.825 ;
        RECT 716.625 50.545 716.905 50.825 ;
        RECT 680.515 50.215 680.795 50.495 ;
        RECT 4.660 47.855 4.940 48.135 ;
        RECT 4.660 47.195 4.940 47.475 ;
        RECT 4.660 46.535 4.940 46.815 ;
        RECT 53.630 45.155 53.910 45.435 ;
        RECT 53.630 44.495 53.910 44.775 ;
        RECT 53.630 43.835 53.910 44.115 ;
        RECT 72.940 42.455 73.220 42.735 ;
        RECT 72.940 41.795 73.220 42.075 ;
        RECT 72.940 41.135 73.220 41.415 ;
        RECT 121.910 39.755 122.190 40.035 ;
        RECT 121.910 39.095 122.190 39.375 ;
        RECT 121.910 38.435 122.190 38.715 ;
        RECT 107.080 30.355 107.360 30.635 ;
        RECT 107.080 29.695 107.360 29.975 ;
        RECT 107.080 29.035 107.360 29.315 ;
        RECT 87.770 27.655 88.050 27.935 ;
        RECT 87.770 26.995 88.050 27.275 ;
        RECT 87.770 26.335 88.050 26.615 ;
        RECT 38.800 24.955 39.080 25.235 ;
        RECT 38.800 24.295 39.080 24.575 ;
        RECT 38.800 23.635 39.080 23.915 ;
        RECT 22.850 22.255 23.130 22.535 ;
        RECT 22.850 21.595 23.130 21.875 ;
        RECT 22.850 20.935 23.130 21.215 ;
        RECT 682.360 18.165 682.640 18.445 ;
        RECT 684.145 18.165 684.425 18.445 ;
        RECT 687.000 18.165 687.280 18.445 ;
        RECT 688.785 18.165 689.065 18.445 ;
        RECT 691.640 18.165 691.920 18.445 ;
        RECT 693.425 18.165 693.705 18.445 ;
        RECT 696.280 18.165 696.560 18.445 ;
        RECT 698.065 18.165 698.345 18.445 ;
        RECT 700.920 18.165 701.200 18.445 ;
        RECT 702.705 18.165 702.985 18.445 ;
        RECT 705.560 18.165 705.840 18.445 ;
        RECT 707.345 18.165 707.625 18.445 ;
        RECT 710.200 18.165 710.480 18.445 ;
        RECT 711.985 18.165 712.265 18.445 ;
        RECT 714.840 18.165 715.120 18.445 ;
        RECT 716.625 18.165 716.905 18.445 ;
        RECT 682.360 17.505 682.640 17.785 ;
        RECT 684.145 17.505 684.425 17.785 ;
        RECT 687.000 17.505 687.280 17.785 ;
        RECT 688.785 17.505 689.065 17.785 ;
        RECT 691.640 17.505 691.920 17.785 ;
        RECT 693.425 17.505 693.705 17.785 ;
        RECT 696.280 17.505 696.560 17.785 ;
        RECT 698.065 17.505 698.345 17.785 ;
        RECT 700.920 17.505 701.200 17.785 ;
        RECT 702.705 17.505 702.985 17.785 ;
        RECT 705.560 17.505 705.840 17.785 ;
        RECT 707.345 17.505 707.625 17.785 ;
        RECT 710.200 17.505 710.480 17.785 ;
        RECT 711.985 17.505 712.265 17.785 ;
        RECT 714.840 17.505 715.120 17.785 ;
        RECT 716.625 17.505 716.905 17.785 ;
        RECT 682.360 16.845 682.640 17.125 ;
        RECT 684.145 16.845 684.425 17.125 ;
        RECT 687.000 16.845 687.280 17.125 ;
        RECT 688.785 16.845 689.065 17.125 ;
        RECT 691.640 16.845 691.920 17.125 ;
        RECT 693.425 16.845 693.705 17.125 ;
        RECT 696.280 16.845 696.560 17.125 ;
        RECT 698.065 16.845 698.345 17.125 ;
        RECT 700.920 16.845 701.200 17.125 ;
        RECT 702.705 16.845 702.985 17.125 ;
        RECT 705.560 16.845 705.840 17.125 ;
        RECT 707.345 16.845 707.625 17.125 ;
        RECT 710.200 16.845 710.480 17.125 ;
        RECT 711.985 16.845 712.265 17.125 ;
        RECT 714.840 16.845 715.120 17.125 ;
        RECT 716.625 16.845 716.905 17.125 ;
        RECT 682.360 16.185 682.640 16.465 ;
        RECT 684.145 16.185 684.425 16.465 ;
        RECT 687.000 16.185 687.280 16.465 ;
        RECT 688.785 16.185 689.065 16.465 ;
        RECT 691.640 16.185 691.920 16.465 ;
        RECT 693.425 16.185 693.705 16.465 ;
        RECT 696.280 16.185 696.560 16.465 ;
        RECT 698.065 16.185 698.345 16.465 ;
        RECT 700.920 16.185 701.200 16.465 ;
        RECT 702.705 16.185 702.985 16.465 ;
        RECT 705.560 16.185 705.840 16.465 ;
        RECT 707.345 16.185 707.625 16.465 ;
        RECT 710.200 16.185 710.480 16.465 ;
        RECT 711.985 16.185 712.265 16.465 ;
        RECT 714.840 16.185 715.120 16.465 ;
        RECT 716.625 16.185 716.905 16.465 ;
        RECT 682.360 15.525 682.640 15.805 ;
        RECT 684.145 15.525 684.425 15.805 ;
        RECT 687.000 15.525 687.280 15.805 ;
        RECT 688.785 15.525 689.065 15.805 ;
        RECT 691.640 15.525 691.920 15.805 ;
        RECT 693.425 15.525 693.705 15.805 ;
        RECT 696.280 15.525 696.560 15.805 ;
        RECT 698.065 15.525 698.345 15.805 ;
        RECT 700.920 15.525 701.200 15.805 ;
        RECT 702.705 15.525 702.985 15.805 ;
        RECT 705.560 15.525 705.840 15.805 ;
        RECT 707.345 15.525 707.625 15.805 ;
        RECT 710.200 15.525 710.480 15.805 ;
        RECT 711.985 15.525 712.265 15.805 ;
        RECT 714.840 15.525 715.120 15.805 ;
        RECT 716.625 15.525 716.905 15.805 ;
        RECT 682.360 14.865 682.640 15.145 ;
        RECT 684.145 14.865 684.425 15.145 ;
        RECT 687.000 14.865 687.280 15.145 ;
        RECT 688.785 14.865 689.065 15.145 ;
        RECT 691.640 14.865 691.920 15.145 ;
        RECT 693.425 14.865 693.705 15.145 ;
        RECT 696.280 14.865 696.560 15.145 ;
        RECT 698.065 14.865 698.345 15.145 ;
        RECT 700.920 14.865 701.200 15.145 ;
        RECT 702.705 14.865 702.985 15.145 ;
        RECT 705.560 14.865 705.840 15.145 ;
        RECT 707.345 14.865 707.625 15.145 ;
        RECT 710.200 14.865 710.480 15.145 ;
        RECT 711.985 14.865 712.265 15.145 ;
        RECT 714.840 14.865 715.120 15.145 ;
        RECT 716.625 14.865 716.905 15.145 ;
        RECT 682.360 14.205 682.640 14.485 ;
        RECT 684.145 14.205 684.425 14.485 ;
        RECT 687.000 14.205 687.280 14.485 ;
        RECT 688.785 14.205 689.065 14.485 ;
        RECT 691.640 14.205 691.920 14.485 ;
        RECT 693.425 14.205 693.705 14.485 ;
        RECT 696.280 14.205 696.560 14.485 ;
        RECT 698.065 14.205 698.345 14.485 ;
        RECT 700.920 14.205 701.200 14.485 ;
        RECT 702.705 14.205 702.985 14.485 ;
        RECT 705.560 14.205 705.840 14.485 ;
        RECT 707.345 14.205 707.625 14.485 ;
        RECT 710.200 14.205 710.480 14.485 ;
        RECT 711.985 14.205 712.265 14.485 ;
        RECT 714.840 14.205 715.120 14.485 ;
        RECT 716.625 14.205 716.905 14.485 ;
        RECT 682.360 13.545 682.640 13.825 ;
        RECT 684.145 13.545 684.425 13.825 ;
        RECT 687.000 13.545 687.280 13.825 ;
        RECT 688.785 13.545 689.065 13.825 ;
        RECT 691.640 13.545 691.920 13.825 ;
        RECT 693.425 13.545 693.705 13.825 ;
        RECT 696.280 13.545 696.560 13.825 ;
        RECT 698.065 13.545 698.345 13.825 ;
        RECT 700.920 13.545 701.200 13.825 ;
        RECT 702.705 13.545 702.985 13.825 ;
        RECT 705.560 13.545 705.840 13.825 ;
        RECT 707.345 13.545 707.625 13.825 ;
        RECT 710.200 13.545 710.480 13.825 ;
        RECT 711.985 13.545 712.265 13.825 ;
        RECT 714.840 13.545 715.120 13.825 ;
        RECT 716.625 13.545 716.905 13.825 ;
        RECT 682.360 12.885 682.640 13.165 ;
        RECT 684.145 12.885 684.425 13.165 ;
        RECT 687.000 12.885 687.280 13.165 ;
        RECT 688.785 12.885 689.065 13.165 ;
        RECT 691.640 12.885 691.920 13.165 ;
        RECT 693.425 12.885 693.705 13.165 ;
        RECT 696.280 12.885 696.560 13.165 ;
        RECT 698.065 12.885 698.345 13.165 ;
        RECT 700.920 12.885 701.200 13.165 ;
        RECT 702.705 12.885 702.985 13.165 ;
        RECT 705.560 12.885 705.840 13.165 ;
        RECT 707.345 12.885 707.625 13.165 ;
        RECT 710.200 12.885 710.480 13.165 ;
        RECT 711.985 12.885 712.265 13.165 ;
        RECT 714.840 12.885 715.120 13.165 ;
        RECT 716.625 12.885 716.905 13.165 ;
        RECT 682.360 12.225 682.640 12.505 ;
        RECT 684.145 12.225 684.425 12.505 ;
        RECT 687.000 12.225 687.280 12.505 ;
        RECT 688.785 12.225 689.065 12.505 ;
        RECT 691.640 12.225 691.920 12.505 ;
        RECT 693.425 12.225 693.705 12.505 ;
        RECT 696.280 12.225 696.560 12.505 ;
        RECT 698.065 12.225 698.345 12.505 ;
        RECT 700.920 12.225 701.200 12.505 ;
        RECT 702.705 12.225 702.985 12.505 ;
        RECT 705.560 12.225 705.840 12.505 ;
        RECT 707.345 12.225 707.625 12.505 ;
        RECT 710.200 12.225 710.480 12.505 ;
        RECT 711.985 12.225 712.265 12.505 ;
        RECT 714.840 12.225 715.120 12.505 ;
        RECT 716.625 12.225 716.905 12.505 ;
        RECT 682.360 11.565 682.640 11.845 ;
        RECT 684.145 11.565 684.425 11.845 ;
        RECT 687.000 11.565 687.280 11.845 ;
        RECT 688.785 11.565 689.065 11.845 ;
        RECT 691.640 11.565 691.920 11.845 ;
        RECT 693.425 11.565 693.705 11.845 ;
        RECT 696.280 11.565 696.560 11.845 ;
        RECT 698.065 11.565 698.345 11.845 ;
        RECT 700.920 11.565 701.200 11.845 ;
        RECT 702.705 11.565 702.985 11.845 ;
        RECT 705.560 11.565 705.840 11.845 ;
        RECT 707.345 11.565 707.625 11.845 ;
        RECT 710.200 11.565 710.480 11.845 ;
        RECT 711.985 11.565 712.265 11.845 ;
        RECT 714.840 11.565 715.120 11.845 ;
        RECT 716.625 11.565 716.905 11.845 ;
        RECT 682.360 10.905 682.640 11.185 ;
        RECT 684.145 10.905 684.425 11.185 ;
        RECT 687.000 10.905 687.280 11.185 ;
        RECT 688.785 10.905 689.065 11.185 ;
        RECT 691.640 10.905 691.920 11.185 ;
        RECT 693.425 10.905 693.705 11.185 ;
        RECT 696.280 10.905 696.560 11.185 ;
        RECT 698.065 10.905 698.345 11.185 ;
        RECT 700.920 10.905 701.200 11.185 ;
        RECT 702.705 10.905 702.985 11.185 ;
        RECT 705.560 10.905 705.840 11.185 ;
        RECT 707.345 10.905 707.625 11.185 ;
        RECT 710.200 10.905 710.480 11.185 ;
        RECT 711.985 10.905 712.265 11.185 ;
        RECT 714.840 10.905 715.120 11.185 ;
        RECT 716.625 10.905 716.905 11.185 ;
        RECT 682.360 10.245 682.640 10.525 ;
        RECT 684.145 10.245 684.425 10.525 ;
        RECT 687.000 10.245 687.280 10.525 ;
        RECT 688.785 10.245 689.065 10.525 ;
        RECT 691.640 10.245 691.920 10.525 ;
        RECT 693.425 10.245 693.705 10.525 ;
        RECT 696.280 10.245 696.560 10.525 ;
        RECT 698.065 10.245 698.345 10.525 ;
        RECT 700.920 10.245 701.200 10.525 ;
        RECT 702.705 10.245 702.985 10.525 ;
        RECT 705.560 10.245 705.840 10.525 ;
        RECT 707.345 10.245 707.625 10.525 ;
        RECT 710.200 10.245 710.480 10.525 ;
        RECT 711.985 10.245 712.265 10.525 ;
        RECT 714.840 10.245 715.120 10.525 ;
        RECT 716.625 10.245 716.905 10.525 ;
        RECT 682.360 9.585 682.640 9.865 ;
        RECT 684.145 9.585 684.425 9.865 ;
        RECT 687.000 9.585 687.280 9.865 ;
        RECT 688.785 9.585 689.065 9.865 ;
        RECT 691.640 9.585 691.920 9.865 ;
        RECT 693.425 9.585 693.705 9.865 ;
        RECT 696.280 9.585 696.560 9.865 ;
        RECT 698.065 9.585 698.345 9.865 ;
        RECT 700.920 9.585 701.200 9.865 ;
        RECT 702.705 9.585 702.985 9.865 ;
        RECT 705.560 9.585 705.840 9.865 ;
        RECT 707.345 9.585 707.625 9.865 ;
        RECT 710.200 9.585 710.480 9.865 ;
        RECT 711.985 9.585 712.265 9.865 ;
        RECT 714.840 9.585 715.120 9.865 ;
        RECT 716.625 9.585 716.905 9.865 ;
        RECT 682.360 8.925 682.640 9.205 ;
        RECT 684.145 8.925 684.425 9.205 ;
        RECT 687.000 8.925 687.280 9.205 ;
        RECT 688.785 8.925 689.065 9.205 ;
        RECT 691.640 8.925 691.920 9.205 ;
        RECT 693.425 8.925 693.705 9.205 ;
        RECT 696.280 8.925 696.560 9.205 ;
        RECT 698.065 8.925 698.345 9.205 ;
        RECT 700.920 8.925 701.200 9.205 ;
        RECT 702.705 8.925 702.985 9.205 ;
        RECT 705.560 8.925 705.840 9.205 ;
        RECT 707.345 8.925 707.625 9.205 ;
        RECT 710.200 8.925 710.480 9.205 ;
        RECT 711.985 8.925 712.265 9.205 ;
        RECT 714.840 8.925 715.120 9.205 ;
        RECT 716.625 8.925 716.905 9.205 ;
        RECT 4.660 8.140 4.940 8.420 ;
        RECT 22.850 8.140 23.130 8.420 ;
        RECT 38.800 8.140 39.080 8.420 ;
        RECT 53.630 8.140 53.910 8.420 ;
        RECT 72.940 8.140 73.220 8.420 ;
        RECT 87.770 8.140 88.050 8.420 ;
        RECT 107.080 8.140 107.360 8.420 ;
        RECT 121.910 8.140 122.190 8.420 ;
        RECT 4.660 7.480 4.940 7.760 ;
        RECT 22.850 7.480 23.130 7.760 ;
        RECT 38.800 7.480 39.080 7.760 ;
        RECT 53.630 7.480 53.910 7.760 ;
        RECT 72.940 7.480 73.220 7.760 ;
        RECT 87.770 7.480 88.050 7.760 ;
        RECT 107.080 7.480 107.360 7.760 ;
        RECT 121.910 7.480 122.190 7.760 ;
        RECT 4.660 6.820 4.940 7.100 ;
        RECT 22.850 6.820 23.130 7.100 ;
        RECT 38.800 6.820 39.080 7.100 ;
        RECT 53.630 6.820 53.910 7.100 ;
        RECT 72.940 6.820 73.220 7.100 ;
        RECT 87.770 6.820 88.050 7.100 ;
        RECT 107.080 6.820 107.360 7.100 ;
        RECT 121.910 6.820 122.190 7.100 ;
        RECT 0.900 4.740 1.180 5.020 ;
        RECT 2.040 4.740 2.320 5.020 ;
        RECT 8.080 4.770 8.360 5.050 ;
        RECT 8.740 4.770 9.020 5.050 ;
        RECT 9.400 4.770 9.680 5.050 ;
        RECT 14.610 4.740 14.890 5.020 ;
        RECT 15.270 4.740 15.550 5.020 ;
        RECT 15.930 4.740 16.210 5.020 ;
        RECT 17.970 4.740 18.250 5.020 ;
        RECT 18.630 4.740 18.910 5.020 ;
        RECT 19.290 4.740 19.570 5.020 ;
        RECT 26.270 4.770 26.550 5.050 ;
        RECT 26.930 4.770 27.210 5.050 ;
        RECT 27.590 4.770 27.870 5.050 ;
        RECT 32.800 4.740 33.080 5.020 ;
        RECT 33.460 4.740 33.740 5.020 ;
        RECT 34.120 4.740 34.400 5.020 ;
        RECT 36.180 4.740 36.460 5.020 ;
        RECT 42.220 4.770 42.500 5.050 ;
        RECT 42.880 4.770 43.160 5.050 ;
        RECT 43.540 4.770 43.820 5.050 ;
        RECT 48.750 4.740 49.030 5.020 ;
        RECT 49.410 4.740 49.690 5.020 ;
        RECT 50.070 4.740 50.350 5.020 ;
        RECT 57.050 4.770 57.330 5.050 ;
        RECT 57.710 4.770 57.990 5.050 ;
        RECT 58.370 4.770 58.650 5.050 ;
        RECT 63.580 4.740 63.860 5.020 ;
        RECT 64.240 4.740 64.520 5.020 ;
        RECT 64.900 4.740 65.180 5.020 ;
        RECT 66.940 4.740 67.220 5.020 ;
        RECT 67.600 4.740 67.880 5.020 ;
        RECT 68.260 4.740 68.540 5.020 ;
        RECT 70.320 4.740 70.600 5.020 ;
        RECT 76.360 4.770 76.640 5.050 ;
        RECT 77.020 4.770 77.300 5.050 ;
        RECT 77.680 4.770 77.960 5.050 ;
        RECT 82.890 4.740 83.170 5.020 ;
        RECT 83.550 4.740 83.830 5.020 ;
        RECT 84.210 4.740 84.490 5.020 ;
        RECT 91.190 4.770 91.470 5.050 ;
        RECT 91.850 4.770 92.130 5.050 ;
        RECT 92.510 4.770 92.790 5.050 ;
        RECT 97.720 4.740 98.000 5.020 ;
        RECT 98.380 4.740 98.660 5.020 ;
        RECT 99.040 4.740 99.320 5.020 ;
        RECT 101.080 4.740 101.360 5.020 ;
        RECT 101.740 4.740 102.020 5.020 ;
        RECT 102.400 4.740 102.680 5.020 ;
        RECT 104.460 4.740 104.740 5.020 ;
        RECT 110.500 4.770 110.780 5.050 ;
        RECT 111.160 4.770 111.440 5.050 ;
        RECT 111.820 4.770 112.100 5.050 ;
        RECT 117.030 4.740 117.310 5.020 ;
        RECT 117.690 4.740 117.970 5.020 ;
        RECT 118.350 4.740 118.630 5.020 ;
        RECT 125.330 4.770 125.610 5.050 ;
        RECT 125.990 4.770 126.270 5.050 ;
        RECT 126.650 4.770 126.930 5.050 ;
        RECT 131.860 4.740 132.140 5.020 ;
        RECT 132.520 4.740 132.800 5.020 ;
        RECT 133.180 4.740 133.460 5.020 ;
        RECT 135.240 4.740 135.520 5.020 ;
        RECT 136.240 4.740 136.520 5.020 ;
        RECT 136.900 4.740 137.180 5.020 ;
        RECT 137.560 4.740 137.840 5.020 ;
        RECT 138.480 4.740 138.760 5.020 ;
        RECT 139.140 4.740 139.420 5.020 ;
        RECT 139.800 4.740 140.080 5.020 ;
        RECT 140.820 4.740 141.100 5.020 ;
        RECT 141.480 4.740 141.760 5.020 ;
        RECT 142.140 4.740 142.420 5.020 ;
        RECT 144.080 4.740 144.360 5.020 ;
        RECT 144.740 4.740 145.020 5.020 ;
        RECT 145.400 4.740 145.680 5.020 ;
        RECT 146.320 4.740 146.600 5.020 ;
        RECT 146.980 4.740 147.260 5.020 ;
        RECT 147.640 4.740 147.920 5.020 ;
        RECT 148.560 4.740 148.840 5.020 ;
        RECT 149.220 4.740 149.500 5.020 ;
        RECT 149.880 4.740 150.160 5.020 ;
        RECT 150.800 4.740 151.080 5.020 ;
        RECT 151.460 4.740 151.740 5.020 ;
        RECT 152.120 4.740 152.400 5.020 ;
        RECT 153.040 4.740 153.320 5.020 ;
        RECT 153.700 4.740 153.980 5.020 ;
        RECT 154.360 4.740 154.640 5.020 ;
        RECT 155.400 4.740 155.680 5.020 ;
        RECT 156.400 4.740 156.680 5.020 ;
        RECT 157.060 4.740 157.340 5.020 ;
        RECT 157.720 4.740 158.000 5.020 ;
        RECT 158.640 4.740 158.920 5.020 ;
        RECT 159.300 4.740 159.580 5.020 ;
        RECT 159.960 4.740 160.240 5.020 ;
        RECT 160.880 4.740 161.160 5.020 ;
        RECT 161.540 4.740 161.820 5.020 ;
        RECT 162.200 4.740 162.480 5.020 ;
        RECT 163.120 4.740 163.400 5.020 ;
        RECT 163.780 4.740 164.060 5.020 ;
        RECT 164.440 4.740 164.720 5.020 ;
        RECT 165.360 4.740 165.640 5.020 ;
        RECT 166.020 4.740 166.300 5.020 ;
        RECT 166.680 4.740 166.960 5.020 ;
        RECT 167.600 4.740 167.880 5.020 ;
        RECT 168.260 4.740 168.540 5.020 ;
        RECT 168.920 4.740 169.200 5.020 ;
        RECT 169.840 4.740 170.120 5.020 ;
        RECT 170.500 4.740 170.780 5.020 ;
        RECT 171.160 4.740 171.440 5.020 ;
        RECT 172.080 4.740 172.360 5.020 ;
        RECT 172.740 4.740 173.020 5.020 ;
        RECT 173.400 4.740 173.680 5.020 ;
        RECT 174.320 4.740 174.600 5.020 ;
        RECT 174.980 4.740 175.260 5.020 ;
        RECT 175.640 4.740 175.920 5.020 ;
        RECT 176.680 4.740 176.960 5.020 ;
        RECT 177.680 4.740 177.960 5.020 ;
        RECT 178.340 4.740 178.620 5.020 ;
        RECT 179.000 4.740 179.280 5.020 ;
        RECT 179.920 4.740 180.200 5.020 ;
        RECT 180.580 4.740 180.860 5.020 ;
        RECT 181.240 4.740 181.520 5.020 ;
        RECT 182.260 4.740 182.540 5.020 ;
        RECT 182.920 4.740 183.200 5.020 ;
        RECT 183.580 4.740 183.860 5.020 ;
        RECT 185.520 4.740 185.800 5.020 ;
        RECT 186.180 4.740 186.460 5.020 ;
        RECT 186.840 4.740 187.120 5.020 ;
        RECT 187.760 4.740 188.040 5.020 ;
        RECT 188.420 4.740 188.700 5.020 ;
        RECT 189.080 4.740 189.360 5.020 ;
        RECT 190.000 4.740 190.280 5.020 ;
        RECT 190.660 4.740 190.940 5.020 ;
        RECT 191.320 4.740 191.600 5.020 ;
        RECT 192.240 4.740 192.520 5.020 ;
        RECT 192.900 4.740 193.180 5.020 ;
        RECT 193.560 4.740 193.840 5.020 ;
        RECT 194.480 4.740 194.760 5.020 ;
        RECT 195.140 4.740 195.420 5.020 ;
        RECT 195.800 4.740 196.080 5.020 ;
        RECT 196.840 4.740 197.120 5.020 ;
        RECT 197.840 4.740 198.120 5.020 ;
        RECT 198.500 4.740 198.780 5.020 ;
        RECT 199.160 4.740 199.440 5.020 ;
        RECT 200.080 4.740 200.360 5.020 ;
        RECT 200.740 4.740 201.020 5.020 ;
        RECT 201.400 4.740 201.680 5.020 ;
        RECT 202.320 4.740 202.600 5.020 ;
        RECT 202.980 4.740 203.260 5.020 ;
        RECT 203.640 4.740 203.920 5.020 ;
        RECT 204.560 4.740 204.840 5.020 ;
        RECT 205.220 4.740 205.500 5.020 ;
        RECT 205.880 4.740 206.160 5.020 ;
        RECT 206.800 4.740 207.080 5.020 ;
        RECT 207.460 4.740 207.740 5.020 ;
        RECT 208.120 4.740 208.400 5.020 ;
        RECT 209.040 4.740 209.320 5.020 ;
        RECT 209.700 4.740 209.980 5.020 ;
        RECT 210.360 4.740 210.640 5.020 ;
        RECT 211.280 4.740 211.560 5.020 ;
        RECT 211.940 4.740 212.220 5.020 ;
        RECT 212.600 4.740 212.880 5.020 ;
        RECT 213.520 4.740 213.800 5.020 ;
        RECT 214.180 4.740 214.460 5.020 ;
        RECT 214.840 4.740 215.120 5.020 ;
        RECT 215.760 4.740 216.040 5.020 ;
        RECT 216.420 4.740 216.700 5.020 ;
        RECT 217.080 4.740 217.360 5.020 ;
        RECT 218.120 4.740 218.400 5.020 ;
        RECT 219.120 4.740 219.400 5.020 ;
        RECT 219.780 4.740 220.060 5.020 ;
        RECT 220.440 4.740 220.720 5.020 ;
        RECT 221.360 4.740 221.640 5.020 ;
        RECT 222.020 4.740 222.300 5.020 ;
        RECT 222.680 4.740 222.960 5.020 ;
        RECT 223.600 4.740 223.880 5.020 ;
        RECT 224.260 4.740 224.540 5.020 ;
        RECT 224.920 4.740 225.200 5.020 ;
        RECT 225.940 4.740 226.220 5.020 ;
        RECT 226.600 4.740 226.880 5.020 ;
        RECT 227.260 4.740 227.540 5.020 ;
        RECT 229.200 4.740 229.480 5.020 ;
        RECT 229.860 4.740 230.140 5.020 ;
        RECT 230.520 4.740 230.800 5.020 ;
        RECT 231.440 4.740 231.720 5.020 ;
        RECT 232.100 4.740 232.380 5.020 ;
        RECT 232.760 4.740 233.040 5.020 ;
        RECT 233.680 4.740 233.960 5.020 ;
        RECT 234.340 4.740 234.620 5.020 ;
        RECT 235.000 4.740 235.280 5.020 ;
        RECT 235.920 4.740 236.200 5.020 ;
        RECT 236.580 4.740 236.860 5.020 ;
        RECT 237.240 4.740 237.520 5.020 ;
        RECT 238.280 4.740 238.560 5.020 ;
        RECT 239.280 4.740 239.560 5.020 ;
        RECT 239.940 4.740 240.220 5.020 ;
        RECT 240.600 4.740 240.880 5.020 ;
        RECT 241.520 4.740 241.800 5.020 ;
        RECT 242.180 4.740 242.460 5.020 ;
        RECT 242.840 4.740 243.120 5.020 ;
        RECT 243.760 4.740 244.040 5.020 ;
        RECT 244.420 4.740 244.700 5.020 ;
        RECT 245.080 4.740 245.360 5.020 ;
        RECT 246.000 4.740 246.280 5.020 ;
        RECT 246.660 4.740 246.940 5.020 ;
        RECT 247.320 4.740 247.600 5.020 ;
        RECT 248.240 4.740 248.520 5.020 ;
        RECT 248.900 4.740 249.180 5.020 ;
        RECT 249.560 4.740 249.840 5.020 ;
        RECT 250.480 4.740 250.760 5.020 ;
        RECT 251.140 4.740 251.420 5.020 ;
        RECT 251.800 4.740 252.080 5.020 ;
        RECT 252.720 4.740 253.000 5.020 ;
        RECT 253.380 4.740 253.660 5.020 ;
        RECT 254.040 4.740 254.320 5.020 ;
        RECT 254.960 4.740 255.240 5.020 ;
        RECT 255.620 4.740 255.900 5.020 ;
        RECT 256.280 4.740 256.560 5.020 ;
        RECT 257.200 4.740 257.480 5.020 ;
        RECT 257.860 4.740 258.140 5.020 ;
        RECT 258.520 4.740 258.800 5.020 ;
        RECT 259.560 4.740 259.840 5.020 ;
        RECT 260.560 4.740 260.840 5.020 ;
        RECT 261.220 4.740 261.500 5.020 ;
        RECT 261.880 4.740 262.160 5.020 ;
        RECT 262.800 4.740 263.080 5.020 ;
        RECT 263.460 4.740 263.740 5.020 ;
        RECT 264.120 4.740 264.400 5.020 ;
        RECT 265.040 4.740 265.320 5.020 ;
        RECT 265.700 4.740 265.980 5.020 ;
        RECT 266.360 4.740 266.640 5.020 ;
        RECT 267.380 4.740 267.660 5.020 ;
        RECT 268.040 4.740 268.320 5.020 ;
        RECT 268.700 4.740 268.980 5.020 ;
        RECT 270.640 4.740 270.920 5.020 ;
        RECT 271.300 4.740 271.580 5.020 ;
        RECT 271.960 4.740 272.240 5.020 ;
        RECT 272.880 4.740 273.160 5.020 ;
        RECT 273.540 4.740 273.820 5.020 ;
        RECT 274.200 4.740 274.480 5.020 ;
        RECT 275.120 4.740 275.400 5.020 ;
        RECT 275.780 4.740 276.060 5.020 ;
        RECT 276.440 4.740 276.720 5.020 ;
        RECT 277.360 4.740 277.640 5.020 ;
        RECT 278.020 4.740 278.300 5.020 ;
        RECT 278.680 4.740 278.960 5.020 ;
        RECT 279.720 4.740 280.000 5.020 ;
        RECT 280.720 4.740 281.000 5.020 ;
        RECT 281.380 4.740 281.660 5.020 ;
        RECT 282.040 4.740 282.320 5.020 ;
        RECT 282.960 4.740 283.240 5.020 ;
        RECT 283.620 4.740 283.900 5.020 ;
        RECT 284.280 4.740 284.560 5.020 ;
        RECT 285.200 4.740 285.480 5.020 ;
        RECT 285.860 4.740 286.140 5.020 ;
        RECT 286.520 4.740 286.800 5.020 ;
        RECT 287.440 4.740 287.720 5.020 ;
        RECT 288.100 4.740 288.380 5.020 ;
        RECT 288.760 4.740 289.040 5.020 ;
        RECT 289.680 4.740 289.960 5.020 ;
        RECT 290.340 4.740 290.620 5.020 ;
        RECT 291.000 4.740 291.280 5.020 ;
        RECT 291.920 4.740 292.200 5.020 ;
        RECT 292.580 4.740 292.860 5.020 ;
        RECT 293.240 4.740 293.520 5.020 ;
        RECT 294.160 4.740 294.440 5.020 ;
        RECT 294.820 4.740 295.100 5.020 ;
        RECT 295.480 4.740 295.760 5.020 ;
        RECT 296.400 4.740 296.680 5.020 ;
        RECT 297.060 4.740 297.340 5.020 ;
        RECT 297.720 4.740 298.000 5.020 ;
        RECT 298.640 4.740 298.920 5.020 ;
        RECT 299.300 4.740 299.580 5.020 ;
        RECT 299.960 4.740 300.240 5.020 ;
        RECT 301.000 4.740 301.280 5.020 ;
        RECT 302.000 4.740 302.280 5.020 ;
        RECT 302.660 4.740 302.940 5.020 ;
        RECT 303.320 4.740 303.600 5.020 ;
        RECT 304.240 4.740 304.520 5.020 ;
        RECT 304.900 4.740 305.180 5.020 ;
        RECT 305.560 4.740 305.840 5.020 ;
        RECT 306.480 4.740 306.760 5.020 ;
        RECT 307.140 4.740 307.420 5.020 ;
        RECT 307.800 4.740 308.080 5.020 ;
        RECT 308.720 4.740 309.000 5.020 ;
        RECT 309.380 4.740 309.660 5.020 ;
        RECT 310.040 4.740 310.320 5.020 ;
        RECT 311.060 4.740 311.340 5.020 ;
        RECT 311.720 4.740 312.000 5.020 ;
        RECT 312.380 4.740 312.660 5.020 ;
        RECT 314.320 4.740 314.600 5.020 ;
        RECT 314.980 4.740 315.260 5.020 ;
        RECT 315.640 4.740 315.920 5.020 ;
        RECT 316.560 4.740 316.840 5.020 ;
        RECT 317.220 4.740 317.500 5.020 ;
        RECT 317.880 4.740 318.160 5.020 ;
        RECT 318.800 4.740 319.080 5.020 ;
        RECT 319.460 4.740 319.740 5.020 ;
        RECT 320.120 4.740 320.400 5.020 ;
        RECT 321.160 4.740 321.440 5.020 ;
        RECT 322.160 4.740 322.440 5.020 ;
        RECT 322.820 4.740 323.100 5.020 ;
        RECT 323.480 4.740 323.760 5.020 ;
        RECT 324.400 4.740 324.680 5.020 ;
        RECT 325.060 4.740 325.340 5.020 ;
        RECT 325.720 4.740 326.000 5.020 ;
        RECT 326.640 4.740 326.920 5.020 ;
        RECT 327.300 4.740 327.580 5.020 ;
        RECT 327.960 4.740 328.240 5.020 ;
        RECT 328.880 4.740 329.160 5.020 ;
        RECT 329.540 4.740 329.820 5.020 ;
        RECT 330.200 4.740 330.480 5.020 ;
        RECT 331.120 4.740 331.400 5.020 ;
        RECT 331.780 4.740 332.060 5.020 ;
        RECT 332.440 4.740 332.720 5.020 ;
        RECT 333.360 4.740 333.640 5.020 ;
        RECT 334.020 4.740 334.300 5.020 ;
        RECT 334.680 4.740 334.960 5.020 ;
        RECT 335.600 4.740 335.880 5.020 ;
        RECT 336.260 4.740 336.540 5.020 ;
        RECT 336.920 4.740 337.200 5.020 ;
        RECT 337.840 4.740 338.120 5.020 ;
        RECT 338.500 4.740 338.780 5.020 ;
        RECT 339.160 4.740 339.440 5.020 ;
        RECT 340.080 4.740 340.360 5.020 ;
        RECT 340.740 4.740 341.020 5.020 ;
        RECT 341.400 4.740 341.680 5.020 ;
        RECT 342.440 4.740 342.720 5.020 ;
        RECT 343.440 4.740 343.720 5.020 ;
        RECT 344.100 4.740 344.380 5.020 ;
        RECT 344.760 4.740 345.040 5.020 ;
        RECT 345.680 4.740 345.960 5.020 ;
        RECT 346.340 4.740 346.620 5.020 ;
        RECT 347.000 4.740 347.280 5.020 ;
        RECT 347.920 4.740 348.200 5.020 ;
        RECT 348.580 4.740 348.860 5.020 ;
        RECT 349.240 4.740 349.520 5.020 ;
        RECT 350.160 4.740 350.440 5.020 ;
        RECT 350.820 4.740 351.100 5.020 ;
        RECT 351.480 4.740 351.760 5.020 ;
        RECT 352.500 4.740 352.780 5.020 ;
        RECT 353.160 4.740 353.440 5.020 ;
        RECT 353.820 4.740 354.100 5.020 ;
        RECT 355.760 4.740 356.040 5.020 ;
        RECT 356.420 4.740 356.700 5.020 ;
        RECT 357.080 4.740 357.360 5.020 ;
        RECT 358.000 4.740 358.280 5.020 ;
        RECT 358.660 4.740 358.940 5.020 ;
        RECT 359.320 4.740 359.600 5.020 ;
        RECT 360.240 4.740 360.520 5.020 ;
        RECT 360.900 4.740 361.180 5.020 ;
        RECT 361.560 4.740 361.840 5.020 ;
        RECT 362.600 4.740 362.880 5.020 ;
        RECT 363.600 4.740 363.880 5.020 ;
        RECT 364.260 4.740 364.540 5.020 ;
        RECT 364.920 4.740 365.200 5.020 ;
        RECT 365.840 4.740 366.120 5.020 ;
        RECT 366.500 4.740 366.780 5.020 ;
        RECT 367.160 4.740 367.440 5.020 ;
        RECT 368.080 4.740 368.360 5.020 ;
        RECT 368.740 4.740 369.020 5.020 ;
        RECT 369.400 4.740 369.680 5.020 ;
        RECT 370.320 4.740 370.600 5.020 ;
        RECT 370.980 4.740 371.260 5.020 ;
        RECT 371.640 4.740 371.920 5.020 ;
        RECT 372.560 4.740 372.840 5.020 ;
        RECT 373.220 4.740 373.500 5.020 ;
        RECT 373.880 4.740 374.160 5.020 ;
        RECT 374.800 4.740 375.080 5.020 ;
        RECT 375.460 4.740 375.740 5.020 ;
        RECT 376.120 4.740 376.400 5.020 ;
        RECT 377.040 4.740 377.320 5.020 ;
        RECT 377.700 4.740 377.980 5.020 ;
        RECT 378.360 4.740 378.640 5.020 ;
        RECT 379.280 4.740 379.560 5.020 ;
        RECT 379.940 4.740 380.220 5.020 ;
        RECT 380.600 4.740 380.880 5.020 ;
        RECT 381.520 4.740 381.800 5.020 ;
        RECT 382.180 4.740 382.460 5.020 ;
        RECT 382.840 4.740 383.120 5.020 ;
        RECT 383.880 4.740 384.160 5.020 ;
        RECT 384.880 4.740 385.160 5.020 ;
        RECT 385.540 4.740 385.820 5.020 ;
        RECT 386.200 4.740 386.480 5.020 ;
        RECT 387.120 4.740 387.400 5.020 ;
        RECT 387.780 4.740 388.060 5.020 ;
        RECT 388.440 4.740 388.720 5.020 ;
        RECT 389.360 4.740 389.640 5.020 ;
        RECT 390.020 4.740 390.300 5.020 ;
        RECT 390.680 4.740 390.960 5.020 ;
        RECT 391.600 4.740 391.880 5.020 ;
        RECT 392.260 4.740 392.540 5.020 ;
        RECT 392.920 4.740 393.200 5.020 ;
        RECT 393.840 4.740 394.120 5.020 ;
        RECT 394.500 4.740 394.780 5.020 ;
        RECT 395.160 4.740 395.440 5.020 ;
        RECT 396.180 4.740 396.460 5.020 ;
        RECT 396.840 4.740 397.120 5.020 ;
        RECT 397.500 4.740 397.780 5.020 ;
        RECT 399.440 4.740 399.720 5.020 ;
        RECT 400.100 4.740 400.380 5.020 ;
        RECT 400.760 4.740 401.040 5.020 ;
        RECT 401.680 4.740 401.960 5.020 ;
        RECT 402.340 4.740 402.620 5.020 ;
        RECT 403.000 4.740 403.280 5.020 ;
        RECT 404.040 4.740 404.320 5.020 ;
        RECT 405.040 4.740 405.320 5.020 ;
        RECT 405.700 4.740 405.980 5.020 ;
        RECT 406.360 4.740 406.640 5.020 ;
        RECT 407.280 4.740 407.560 5.020 ;
        RECT 407.940 4.740 408.220 5.020 ;
        RECT 408.600 4.740 408.880 5.020 ;
        RECT 409.520 4.740 409.800 5.020 ;
        RECT 410.180 4.740 410.460 5.020 ;
        RECT 410.840 4.740 411.120 5.020 ;
        RECT 411.760 4.740 412.040 5.020 ;
        RECT 412.420 4.740 412.700 5.020 ;
        RECT 413.080 4.740 413.360 5.020 ;
        RECT 414.000 4.740 414.280 5.020 ;
        RECT 414.660 4.740 414.940 5.020 ;
        RECT 415.320 4.740 415.600 5.020 ;
        RECT 416.240 4.740 416.520 5.020 ;
        RECT 416.900 4.740 417.180 5.020 ;
        RECT 417.560 4.740 417.840 5.020 ;
        RECT 418.480 4.740 418.760 5.020 ;
        RECT 419.140 4.740 419.420 5.020 ;
        RECT 419.800 4.740 420.080 5.020 ;
        RECT 420.720 4.740 421.000 5.020 ;
        RECT 421.380 4.740 421.660 5.020 ;
        RECT 422.040 4.740 422.320 5.020 ;
        RECT 422.960 4.740 423.240 5.020 ;
        RECT 423.620 4.740 423.900 5.020 ;
        RECT 424.280 4.740 424.560 5.020 ;
        RECT 425.320 4.740 425.600 5.020 ;
        RECT 426.320 4.740 426.600 5.020 ;
        RECT 426.980 4.740 427.260 5.020 ;
        RECT 427.640 4.740 427.920 5.020 ;
        RECT 428.560 4.740 428.840 5.020 ;
        RECT 429.220 4.740 429.500 5.020 ;
        RECT 429.880 4.740 430.160 5.020 ;
        RECT 430.800 4.740 431.080 5.020 ;
        RECT 431.460 4.740 431.740 5.020 ;
        RECT 432.120 4.740 432.400 5.020 ;
        RECT 433.040 4.740 433.320 5.020 ;
        RECT 433.700 4.740 433.980 5.020 ;
        RECT 434.360 4.740 434.640 5.020 ;
        RECT 435.280 4.740 435.560 5.020 ;
        RECT 435.940 4.740 436.220 5.020 ;
        RECT 436.600 4.740 436.880 5.020 ;
        RECT 437.620 4.740 437.900 5.020 ;
        RECT 438.280 4.740 438.560 5.020 ;
        RECT 438.940 4.740 439.220 5.020 ;
        RECT 440.880 4.740 441.160 5.020 ;
        RECT 441.540 4.740 441.820 5.020 ;
        RECT 442.200 4.740 442.480 5.020 ;
        RECT 443.120 4.740 443.400 5.020 ;
        RECT 443.780 4.740 444.060 5.020 ;
        RECT 444.440 4.740 444.720 5.020 ;
        RECT 445.480 4.740 445.760 5.020 ;
        RECT 446.480 4.740 446.760 5.020 ;
        RECT 447.140 4.740 447.420 5.020 ;
        RECT 447.800 4.740 448.080 5.020 ;
        RECT 448.720 4.740 449.000 5.020 ;
        RECT 449.380 4.740 449.660 5.020 ;
        RECT 450.040 4.740 450.320 5.020 ;
        RECT 450.960 4.740 451.240 5.020 ;
        RECT 451.620 4.740 451.900 5.020 ;
        RECT 452.280 4.740 452.560 5.020 ;
        RECT 453.200 4.740 453.480 5.020 ;
        RECT 453.860 4.740 454.140 5.020 ;
        RECT 454.520 4.740 454.800 5.020 ;
        RECT 455.440 4.740 455.720 5.020 ;
        RECT 456.100 4.740 456.380 5.020 ;
        RECT 456.760 4.740 457.040 5.020 ;
        RECT 457.680 4.740 457.960 5.020 ;
        RECT 458.340 4.740 458.620 5.020 ;
        RECT 459.000 4.740 459.280 5.020 ;
        RECT 459.920 4.740 460.200 5.020 ;
        RECT 460.580 4.740 460.860 5.020 ;
        RECT 461.240 4.740 461.520 5.020 ;
        RECT 462.160 4.740 462.440 5.020 ;
        RECT 462.820 4.740 463.100 5.020 ;
        RECT 463.480 4.740 463.760 5.020 ;
        RECT 464.400 4.740 464.680 5.020 ;
        RECT 465.060 4.740 465.340 5.020 ;
        RECT 465.720 4.740 466.000 5.020 ;
        RECT 466.760 4.740 467.040 5.020 ;
        RECT 467.760 4.740 468.040 5.020 ;
        RECT 468.420 4.740 468.700 5.020 ;
        RECT 469.080 4.740 469.360 5.020 ;
        RECT 470.000 4.740 470.280 5.020 ;
        RECT 470.660 4.740 470.940 5.020 ;
        RECT 471.320 4.740 471.600 5.020 ;
        RECT 472.240 4.740 472.520 5.020 ;
        RECT 472.900 4.740 473.180 5.020 ;
        RECT 473.560 4.740 473.840 5.020 ;
        RECT 474.480 4.740 474.760 5.020 ;
        RECT 475.140 4.740 475.420 5.020 ;
        RECT 475.800 4.740 476.080 5.020 ;
        RECT 476.720 4.740 477.000 5.020 ;
        RECT 477.380 4.740 477.660 5.020 ;
        RECT 478.040 4.740 478.320 5.020 ;
        RECT 478.960 4.740 479.240 5.020 ;
        RECT 479.620 4.740 479.900 5.020 ;
        RECT 480.280 4.740 480.560 5.020 ;
        RECT 481.300 4.740 481.580 5.020 ;
        RECT 481.960 4.740 482.240 5.020 ;
        RECT 482.620 4.740 482.900 5.020 ;
        RECT 484.560 4.740 484.840 5.020 ;
        RECT 485.220 4.740 485.500 5.020 ;
        RECT 485.880 4.740 486.160 5.020 ;
        RECT 486.920 4.740 487.200 5.020 ;
        RECT 487.920 4.740 488.200 5.020 ;
        RECT 488.580 4.740 488.860 5.020 ;
        RECT 489.240 4.740 489.520 5.020 ;
        RECT 490.160 4.740 490.440 5.020 ;
        RECT 490.820 4.740 491.100 5.020 ;
        RECT 491.480 4.740 491.760 5.020 ;
        RECT 492.400 4.740 492.680 5.020 ;
        RECT 493.060 4.740 493.340 5.020 ;
        RECT 493.720 4.740 494.000 5.020 ;
        RECT 494.640 4.740 494.920 5.020 ;
        RECT 495.300 4.740 495.580 5.020 ;
        RECT 495.960 4.740 496.240 5.020 ;
        RECT 496.880 4.740 497.160 5.020 ;
        RECT 497.540 4.740 497.820 5.020 ;
        RECT 498.200 4.740 498.480 5.020 ;
        RECT 499.120 4.740 499.400 5.020 ;
        RECT 499.780 4.740 500.060 5.020 ;
        RECT 500.440 4.740 500.720 5.020 ;
        RECT 501.360 4.740 501.640 5.020 ;
        RECT 502.020 4.740 502.300 5.020 ;
        RECT 502.680 4.740 502.960 5.020 ;
        RECT 503.600 4.740 503.880 5.020 ;
        RECT 504.260 4.740 504.540 5.020 ;
        RECT 504.920 4.740 505.200 5.020 ;
        RECT 505.840 4.740 506.120 5.020 ;
        RECT 506.500 4.740 506.780 5.020 ;
        RECT 507.160 4.740 507.440 5.020 ;
        RECT 508.200 4.740 508.480 5.020 ;
        RECT 509.200 4.740 509.480 5.020 ;
        RECT 509.860 4.740 510.140 5.020 ;
        RECT 510.520 4.740 510.800 5.020 ;
        RECT 511.440 4.740 511.720 5.020 ;
        RECT 512.100 4.740 512.380 5.020 ;
        RECT 512.760 4.740 513.040 5.020 ;
        RECT 513.680 4.740 513.960 5.020 ;
        RECT 514.340 4.740 514.620 5.020 ;
        RECT 515.000 4.740 515.280 5.020 ;
        RECT 515.920 4.740 516.200 5.020 ;
        RECT 516.580 4.740 516.860 5.020 ;
        RECT 517.240 4.740 517.520 5.020 ;
        RECT 518.160 4.740 518.440 5.020 ;
        RECT 518.820 4.740 519.100 5.020 ;
        RECT 519.480 4.740 519.760 5.020 ;
        RECT 520.400 4.740 520.680 5.020 ;
        RECT 521.060 4.740 521.340 5.020 ;
        RECT 521.720 4.740 522.000 5.020 ;
        RECT 522.740 4.740 523.020 5.020 ;
        RECT 523.400 4.740 523.680 5.020 ;
        RECT 524.060 4.740 524.340 5.020 ;
        RECT 526.000 4.740 526.280 5.020 ;
        RECT 526.660 4.740 526.940 5.020 ;
        RECT 527.320 4.740 527.600 5.020 ;
        RECT 528.360 4.740 528.640 5.020 ;
        RECT 529.360 4.740 529.640 5.020 ;
        RECT 530.020 4.740 530.300 5.020 ;
        RECT 530.680 4.740 530.960 5.020 ;
        RECT 531.600 4.740 531.880 5.020 ;
        RECT 532.260 4.740 532.540 5.020 ;
        RECT 532.920 4.740 533.200 5.020 ;
        RECT 533.840 4.740 534.120 5.020 ;
        RECT 534.500 4.740 534.780 5.020 ;
        RECT 535.160 4.740 535.440 5.020 ;
        RECT 536.080 4.740 536.360 5.020 ;
        RECT 536.740 4.740 537.020 5.020 ;
        RECT 537.400 4.740 537.680 5.020 ;
        RECT 538.320 4.740 538.600 5.020 ;
        RECT 538.980 4.740 539.260 5.020 ;
        RECT 539.640 4.740 539.920 5.020 ;
        RECT 540.560 4.740 540.840 5.020 ;
        RECT 541.220 4.740 541.500 5.020 ;
        RECT 541.880 4.740 542.160 5.020 ;
        RECT 542.800 4.740 543.080 5.020 ;
        RECT 543.460 4.740 543.740 5.020 ;
        RECT 544.120 4.740 544.400 5.020 ;
        RECT 545.040 4.740 545.320 5.020 ;
        RECT 545.700 4.740 545.980 5.020 ;
        RECT 546.360 4.740 546.640 5.020 ;
        RECT 547.280 4.740 547.560 5.020 ;
        RECT 547.940 4.740 548.220 5.020 ;
        RECT 548.600 4.740 548.880 5.020 ;
        RECT 549.640 4.740 549.920 5.020 ;
        RECT 550.640 4.740 550.920 5.020 ;
        RECT 551.300 4.740 551.580 5.020 ;
        RECT 551.960 4.740 552.240 5.020 ;
        RECT 552.880 4.740 553.160 5.020 ;
        RECT 553.540 4.740 553.820 5.020 ;
        RECT 554.200 4.740 554.480 5.020 ;
        RECT 555.120 4.740 555.400 5.020 ;
        RECT 555.780 4.740 556.060 5.020 ;
        RECT 556.440 4.740 556.720 5.020 ;
        RECT 557.360 4.740 557.640 5.020 ;
        RECT 558.020 4.740 558.300 5.020 ;
        RECT 558.680 4.740 558.960 5.020 ;
        RECT 559.600 4.740 559.880 5.020 ;
        RECT 560.260 4.740 560.540 5.020 ;
        RECT 560.920 4.740 561.200 5.020 ;
        RECT 561.840 4.740 562.120 5.020 ;
        RECT 562.500 4.740 562.780 5.020 ;
        RECT 563.160 4.740 563.440 5.020 ;
        RECT 564.080 4.740 564.360 5.020 ;
        RECT 564.740 4.740 565.020 5.020 ;
        RECT 565.400 4.740 565.680 5.020 ;
        RECT 566.420 4.740 566.700 5.020 ;
        RECT 567.080 4.740 567.360 5.020 ;
        RECT 567.740 4.740 568.020 5.020 ;
        RECT 569.800 4.740 570.080 5.020 ;
        RECT 570.800 4.740 571.080 5.020 ;
        RECT 571.460 4.740 571.740 5.020 ;
        RECT 572.120 4.740 572.400 5.020 ;
        RECT 573.040 4.740 573.320 5.020 ;
        RECT 573.700 4.740 573.980 5.020 ;
        RECT 574.360 4.740 574.640 5.020 ;
        RECT 575.280 4.740 575.560 5.020 ;
        RECT 575.940 4.740 576.220 5.020 ;
        RECT 576.600 4.740 576.880 5.020 ;
        RECT 577.520 4.740 577.800 5.020 ;
        RECT 578.180 4.740 578.460 5.020 ;
        RECT 578.840 4.740 579.120 5.020 ;
        RECT 579.760 4.740 580.040 5.020 ;
        RECT 580.420 4.740 580.700 5.020 ;
        RECT 581.080 4.740 581.360 5.020 ;
        RECT 582.000 4.740 582.280 5.020 ;
        RECT 582.660 4.740 582.940 5.020 ;
        RECT 583.320 4.740 583.600 5.020 ;
        RECT 584.240 4.740 584.520 5.020 ;
        RECT 584.900 4.740 585.180 5.020 ;
        RECT 585.560 4.740 585.840 5.020 ;
        RECT 586.480 4.740 586.760 5.020 ;
        RECT 587.140 4.740 587.420 5.020 ;
        RECT 587.800 4.740 588.080 5.020 ;
        RECT 588.720 4.740 589.000 5.020 ;
        RECT 589.380 4.740 589.660 5.020 ;
        RECT 590.040 4.740 590.320 5.020 ;
        RECT 591.080 4.740 591.360 5.020 ;
        RECT 592.080 4.740 592.360 5.020 ;
        RECT 592.740 4.740 593.020 5.020 ;
        RECT 593.400 4.740 593.680 5.020 ;
        RECT 594.320 4.740 594.600 5.020 ;
        RECT 594.980 4.740 595.260 5.020 ;
        RECT 595.640 4.740 595.920 5.020 ;
        RECT 596.560 4.740 596.840 5.020 ;
        RECT 597.220 4.740 597.500 5.020 ;
        RECT 597.880 4.740 598.160 5.020 ;
        RECT 598.800 4.740 599.080 5.020 ;
        RECT 599.460 4.740 599.740 5.020 ;
        RECT 600.120 4.740 600.400 5.020 ;
        RECT 601.040 4.740 601.320 5.020 ;
        RECT 601.700 4.740 601.980 5.020 ;
        RECT 602.360 4.740 602.640 5.020 ;
        RECT 603.280 4.740 603.560 5.020 ;
        RECT 603.940 4.740 604.220 5.020 ;
        RECT 604.600 4.740 604.880 5.020 ;
        RECT 605.520 4.740 605.800 5.020 ;
        RECT 606.180 4.740 606.460 5.020 ;
        RECT 606.840 4.740 607.120 5.020 ;
        RECT 607.860 4.740 608.140 5.020 ;
        RECT 608.520 4.740 608.800 5.020 ;
        RECT 609.180 4.740 609.460 5.020 ;
        RECT 611.240 4.740 611.520 5.020 ;
        RECT 612.240 4.740 612.520 5.020 ;
        RECT 612.900 4.740 613.180 5.020 ;
        RECT 613.560 4.740 613.840 5.020 ;
        RECT 614.480 4.740 614.760 5.020 ;
        RECT 615.140 4.740 615.420 5.020 ;
        RECT 615.800 4.740 616.080 5.020 ;
        RECT 616.720 4.740 617.000 5.020 ;
        RECT 617.380 4.740 617.660 5.020 ;
        RECT 618.040 4.740 618.320 5.020 ;
        RECT 618.960 4.740 619.240 5.020 ;
        RECT 619.620 4.740 619.900 5.020 ;
        RECT 620.280 4.740 620.560 5.020 ;
        RECT 621.200 4.740 621.480 5.020 ;
        RECT 621.860 4.740 622.140 5.020 ;
        RECT 622.520 4.740 622.800 5.020 ;
        RECT 623.440 4.740 623.720 5.020 ;
        RECT 624.100 4.740 624.380 5.020 ;
        RECT 624.760 4.740 625.040 5.020 ;
        RECT 625.680 4.740 625.960 5.020 ;
        RECT 626.340 4.740 626.620 5.020 ;
        RECT 627.000 4.740 627.280 5.020 ;
        RECT 627.920 4.740 628.200 5.020 ;
        RECT 628.580 4.740 628.860 5.020 ;
        RECT 629.240 4.740 629.520 5.020 ;
        RECT 630.160 4.740 630.440 5.020 ;
        RECT 630.820 4.740 631.100 5.020 ;
        RECT 631.480 4.740 631.760 5.020 ;
        RECT 632.520 4.740 632.800 5.020 ;
        RECT 633.520 4.740 633.800 5.020 ;
        RECT 634.180 4.740 634.460 5.020 ;
        RECT 634.840 4.740 635.120 5.020 ;
        RECT 635.760 4.740 636.040 5.020 ;
        RECT 636.420 4.740 636.700 5.020 ;
        RECT 637.080 4.740 637.360 5.020 ;
        RECT 638.000 4.740 638.280 5.020 ;
        RECT 638.660 4.740 638.940 5.020 ;
        RECT 639.320 4.740 639.600 5.020 ;
        RECT 640.240 4.740 640.520 5.020 ;
        RECT 640.900 4.740 641.180 5.020 ;
        RECT 641.560 4.740 641.840 5.020 ;
        RECT 642.480 4.740 642.760 5.020 ;
        RECT 643.140 4.740 643.420 5.020 ;
        RECT 643.800 4.740 644.080 5.020 ;
        RECT 644.720 4.740 645.000 5.020 ;
        RECT 645.380 4.740 645.660 5.020 ;
        RECT 646.040 4.740 646.320 5.020 ;
        RECT 646.960 4.740 647.240 5.020 ;
        RECT 647.620 4.740 647.900 5.020 ;
        RECT 648.280 4.740 648.560 5.020 ;
        RECT 649.200 4.740 649.480 5.020 ;
        RECT 649.860 4.740 650.140 5.020 ;
        RECT 650.520 4.740 650.800 5.020 ;
        RECT 651.540 4.740 651.820 5.020 ;
        RECT 652.200 4.740 652.480 5.020 ;
        RECT 652.860 4.740 653.140 5.020 ;
        RECT 654.920 4.740 655.200 5.020 ;
        RECT 655.920 4.740 656.200 5.020 ;
        RECT 656.580 4.740 656.860 5.020 ;
        RECT 657.240 4.740 657.520 5.020 ;
        RECT 658.160 4.740 658.440 5.020 ;
        RECT 658.820 4.740 659.100 5.020 ;
        RECT 659.480 4.740 659.760 5.020 ;
        RECT 660.400 4.740 660.680 5.020 ;
        RECT 661.060 4.740 661.340 5.020 ;
        RECT 661.720 4.740 662.000 5.020 ;
        RECT 662.640 4.740 662.920 5.020 ;
        RECT 663.300 4.740 663.580 5.020 ;
        RECT 663.960 4.740 664.240 5.020 ;
        RECT 664.880 4.740 665.160 5.020 ;
        RECT 665.540 4.740 665.820 5.020 ;
        RECT 666.200 4.740 666.480 5.020 ;
        RECT 667.120 4.740 667.400 5.020 ;
        RECT 667.780 4.740 668.060 5.020 ;
        RECT 668.440 4.740 668.720 5.020 ;
        RECT 669.360 4.740 669.640 5.020 ;
        RECT 670.020 4.740 670.300 5.020 ;
        RECT 670.680 4.740 670.960 5.020 ;
        RECT 671.600 4.740 671.880 5.020 ;
        RECT 672.260 4.740 672.540 5.020 ;
        RECT 672.920 4.740 673.200 5.020 ;
        RECT 673.840 4.740 674.120 5.020 ;
        RECT 674.500 4.740 674.780 5.020 ;
        RECT 675.160 4.740 675.440 5.020 ;
        RECT 676.200 4.740 676.480 5.020 ;
        RECT 677.200 4.740 677.480 5.020 ;
        RECT 677.860 4.740 678.140 5.020 ;
        RECT 678.520 4.740 678.800 5.020 ;
        RECT 679.540 4.740 679.820 5.020 ;
        RECT 0.900 0.820 1.180 1.100 ;
        RECT 2.040 0.820 2.320 1.100 ;
        RECT 7.480 0.820 7.760 1.100 ;
        RECT 8.140 0.820 8.420 1.100 ;
        RECT 8.800 0.820 9.080 1.100 ;
        RECT 14.350 0.820 14.630 1.100 ;
        RECT 15.670 0.820 15.950 1.100 ;
        RECT 17.710 0.820 17.990 1.100 ;
        RECT 19.030 0.820 19.310 1.100 ;
        RECT 25.670 0.820 25.950 1.100 ;
        RECT 26.330 0.820 26.610 1.100 ;
        RECT 26.990 0.820 27.270 1.100 ;
        RECT 32.540 0.820 32.820 1.100 ;
        RECT 33.860 0.820 34.140 1.100 ;
        RECT 36.180 0.820 36.460 1.100 ;
        RECT 41.620 0.820 41.900 1.100 ;
        RECT 42.280 0.820 42.560 1.100 ;
        RECT 42.940 0.820 43.220 1.100 ;
        RECT 48.490 0.820 48.770 1.100 ;
        RECT 49.810 0.820 50.090 1.100 ;
        RECT 56.450 0.820 56.730 1.100 ;
        RECT 57.110 0.820 57.390 1.100 ;
        RECT 57.770 0.820 58.050 1.100 ;
        RECT 63.320 0.820 63.600 1.100 ;
        RECT 64.640 0.820 64.920 1.100 ;
        RECT 66.680 0.820 66.960 1.100 ;
        RECT 68.000 0.820 68.280 1.100 ;
        RECT 70.320 0.820 70.600 1.100 ;
        RECT 75.760 0.820 76.040 1.100 ;
        RECT 76.420 0.820 76.700 1.100 ;
        RECT 77.080 0.820 77.360 1.100 ;
        RECT 82.630 0.820 82.910 1.100 ;
        RECT 83.950 0.820 84.230 1.100 ;
        RECT 90.590 0.820 90.870 1.100 ;
        RECT 91.250 0.820 91.530 1.100 ;
        RECT 91.910 0.820 92.190 1.100 ;
        RECT 97.460 0.820 97.740 1.100 ;
        RECT 98.780 0.820 99.060 1.100 ;
        RECT 100.820 0.820 101.100 1.100 ;
        RECT 102.140 0.820 102.420 1.100 ;
        RECT 104.460 0.820 104.740 1.100 ;
        RECT 109.900 0.820 110.180 1.100 ;
        RECT 110.560 0.820 110.840 1.100 ;
        RECT 111.220 0.820 111.500 1.100 ;
        RECT 116.770 0.820 117.050 1.100 ;
        RECT 118.090 0.820 118.370 1.100 ;
        RECT 124.730 0.820 125.010 1.100 ;
        RECT 125.390 0.820 125.670 1.100 ;
        RECT 126.050 0.820 126.330 1.100 ;
        RECT 131.600 0.820 131.880 1.100 ;
        RECT 132.920 0.820 133.200 1.100 ;
        RECT 135.240 0.820 135.520 1.100 ;
        RECT 136.240 0.820 136.520 1.100 ;
        RECT 136.900 0.820 137.180 1.100 ;
        RECT 137.560 0.820 137.840 1.100 ;
        RECT 138.480 0.820 138.760 1.100 ;
        RECT 139.140 0.820 139.420 1.100 ;
        RECT 139.800 0.820 140.080 1.100 ;
        RECT 140.560 0.820 140.840 1.100 ;
        RECT 141.880 0.820 142.160 1.100 ;
        RECT 144.080 0.820 144.360 1.100 ;
        RECT 144.740 0.820 145.020 1.100 ;
        RECT 145.400 0.820 145.680 1.100 ;
        RECT 146.320 0.820 146.600 1.100 ;
        RECT 146.980 0.820 147.260 1.100 ;
        RECT 147.640 0.820 147.920 1.100 ;
        RECT 148.560 0.820 148.840 1.100 ;
        RECT 149.220 0.820 149.500 1.100 ;
        RECT 149.880 0.820 150.160 1.100 ;
        RECT 150.800 0.820 151.080 1.100 ;
        RECT 151.460 0.820 151.740 1.100 ;
        RECT 152.120 0.820 152.400 1.100 ;
        RECT 153.040 0.820 153.320 1.100 ;
        RECT 153.700 0.820 153.980 1.100 ;
        RECT 154.360 0.820 154.640 1.100 ;
        RECT 155.400 0.820 155.680 1.100 ;
        RECT 156.400 0.820 156.680 1.100 ;
        RECT 157.060 0.820 157.340 1.100 ;
        RECT 157.720 0.820 158.000 1.100 ;
        RECT 158.640 0.820 158.920 1.100 ;
        RECT 159.300 0.820 159.580 1.100 ;
        RECT 159.960 0.820 160.240 1.100 ;
        RECT 160.880 0.820 161.160 1.100 ;
        RECT 161.540 0.820 161.820 1.100 ;
        RECT 162.200 0.820 162.480 1.100 ;
        RECT 163.120 0.820 163.400 1.100 ;
        RECT 163.780 0.820 164.060 1.100 ;
        RECT 164.440 0.820 164.720 1.100 ;
        RECT 165.360 0.820 165.640 1.100 ;
        RECT 166.020 0.820 166.300 1.100 ;
        RECT 166.680 0.820 166.960 1.100 ;
        RECT 167.600 0.820 167.880 1.100 ;
        RECT 168.260 0.820 168.540 1.100 ;
        RECT 168.920 0.820 169.200 1.100 ;
        RECT 169.840 0.820 170.120 1.100 ;
        RECT 170.500 0.820 170.780 1.100 ;
        RECT 171.160 0.820 171.440 1.100 ;
        RECT 172.080 0.820 172.360 1.100 ;
        RECT 172.740 0.820 173.020 1.100 ;
        RECT 173.400 0.820 173.680 1.100 ;
        RECT 174.320 0.820 174.600 1.100 ;
        RECT 174.980 0.820 175.260 1.100 ;
        RECT 175.640 0.820 175.920 1.100 ;
        RECT 176.680 0.820 176.960 1.100 ;
        RECT 177.680 0.820 177.960 1.100 ;
        RECT 178.340 0.820 178.620 1.100 ;
        RECT 179.000 0.820 179.280 1.100 ;
        RECT 179.920 0.820 180.200 1.100 ;
        RECT 180.580 0.820 180.860 1.100 ;
        RECT 181.240 0.820 181.520 1.100 ;
        RECT 182.000 0.820 182.280 1.100 ;
        RECT 183.320 0.820 183.600 1.100 ;
        RECT 185.520 0.820 185.800 1.100 ;
        RECT 186.180 0.820 186.460 1.100 ;
        RECT 186.840 0.820 187.120 1.100 ;
        RECT 187.760 0.820 188.040 1.100 ;
        RECT 188.420 0.820 188.700 1.100 ;
        RECT 189.080 0.820 189.360 1.100 ;
        RECT 190.000 0.820 190.280 1.100 ;
        RECT 190.660 0.820 190.940 1.100 ;
        RECT 191.320 0.820 191.600 1.100 ;
        RECT 192.240 0.820 192.520 1.100 ;
        RECT 192.900 0.820 193.180 1.100 ;
        RECT 193.560 0.820 193.840 1.100 ;
        RECT 194.480 0.820 194.760 1.100 ;
        RECT 195.140 0.820 195.420 1.100 ;
        RECT 195.800 0.820 196.080 1.100 ;
        RECT 196.840 0.820 197.120 1.100 ;
        RECT 197.840 0.820 198.120 1.100 ;
        RECT 198.500 0.820 198.780 1.100 ;
        RECT 199.160 0.820 199.440 1.100 ;
        RECT 200.080 0.820 200.360 1.100 ;
        RECT 200.740 0.820 201.020 1.100 ;
        RECT 201.400 0.820 201.680 1.100 ;
        RECT 202.320 0.820 202.600 1.100 ;
        RECT 202.980 0.820 203.260 1.100 ;
        RECT 203.640 0.820 203.920 1.100 ;
        RECT 204.560 0.820 204.840 1.100 ;
        RECT 205.220 0.820 205.500 1.100 ;
        RECT 205.880 0.820 206.160 1.100 ;
        RECT 206.800 0.820 207.080 1.100 ;
        RECT 207.460 0.820 207.740 1.100 ;
        RECT 208.120 0.820 208.400 1.100 ;
        RECT 209.040 0.820 209.320 1.100 ;
        RECT 209.700 0.820 209.980 1.100 ;
        RECT 210.360 0.820 210.640 1.100 ;
        RECT 211.280 0.820 211.560 1.100 ;
        RECT 211.940 0.820 212.220 1.100 ;
        RECT 212.600 0.820 212.880 1.100 ;
        RECT 213.520 0.820 213.800 1.100 ;
        RECT 214.180 0.820 214.460 1.100 ;
        RECT 214.840 0.820 215.120 1.100 ;
        RECT 215.760 0.820 216.040 1.100 ;
        RECT 216.420 0.820 216.700 1.100 ;
        RECT 217.080 0.820 217.360 1.100 ;
        RECT 218.120 0.820 218.400 1.100 ;
        RECT 219.120 0.820 219.400 1.100 ;
        RECT 219.780 0.820 220.060 1.100 ;
        RECT 220.440 0.820 220.720 1.100 ;
        RECT 221.360 0.820 221.640 1.100 ;
        RECT 222.020 0.820 222.300 1.100 ;
        RECT 222.680 0.820 222.960 1.100 ;
        RECT 223.600 0.820 223.880 1.100 ;
        RECT 224.260 0.820 224.540 1.100 ;
        RECT 224.920 0.820 225.200 1.100 ;
        RECT 225.680 0.820 225.960 1.100 ;
        RECT 227.000 0.820 227.280 1.100 ;
        RECT 229.200 0.820 229.480 1.100 ;
        RECT 229.860 0.820 230.140 1.100 ;
        RECT 230.520 0.820 230.800 1.100 ;
        RECT 231.440 0.820 231.720 1.100 ;
        RECT 232.100 0.820 232.380 1.100 ;
        RECT 232.760 0.820 233.040 1.100 ;
        RECT 233.680 0.820 233.960 1.100 ;
        RECT 234.340 0.820 234.620 1.100 ;
        RECT 235.000 0.820 235.280 1.100 ;
        RECT 235.920 0.820 236.200 1.100 ;
        RECT 236.580 0.820 236.860 1.100 ;
        RECT 237.240 0.820 237.520 1.100 ;
        RECT 238.280 0.820 238.560 1.100 ;
        RECT 239.280 0.820 239.560 1.100 ;
        RECT 239.940 0.820 240.220 1.100 ;
        RECT 240.600 0.820 240.880 1.100 ;
        RECT 241.520 0.820 241.800 1.100 ;
        RECT 242.180 0.820 242.460 1.100 ;
        RECT 242.840 0.820 243.120 1.100 ;
        RECT 243.760 0.820 244.040 1.100 ;
        RECT 244.420 0.820 244.700 1.100 ;
        RECT 245.080 0.820 245.360 1.100 ;
        RECT 246.000 0.820 246.280 1.100 ;
        RECT 246.660 0.820 246.940 1.100 ;
        RECT 247.320 0.820 247.600 1.100 ;
        RECT 248.240 0.820 248.520 1.100 ;
        RECT 248.900 0.820 249.180 1.100 ;
        RECT 249.560 0.820 249.840 1.100 ;
        RECT 250.480 0.820 250.760 1.100 ;
        RECT 251.140 0.820 251.420 1.100 ;
        RECT 251.800 0.820 252.080 1.100 ;
        RECT 252.720 0.820 253.000 1.100 ;
        RECT 253.380 0.820 253.660 1.100 ;
        RECT 254.040 0.820 254.320 1.100 ;
        RECT 254.960 0.820 255.240 1.100 ;
        RECT 255.620 0.820 255.900 1.100 ;
        RECT 256.280 0.820 256.560 1.100 ;
        RECT 257.200 0.820 257.480 1.100 ;
        RECT 257.860 0.820 258.140 1.100 ;
        RECT 258.520 0.820 258.800 1.100 ;
        RECT 259.560 0.820 259.840 1.100 ;
        RECT 260.560 0.820 260.840 1.100 ;
        RECT 261.220 0.820 261.500 1.100 ;
        RECT 261.880 0.820 262.160 1.100 ;
        RECT 262.800 0.820 263.080 1.100 ;
        RECT 263.460 0.820 263.740 1.100 ;
        RECT 264.120 0.820 264.400 1.100 ;
        RECT 265.040 0.820 265.320 1.100 ;
        RECT 265.700 0.820 265.980 1.100 ;
        RECT 266.360 0.820 266.640 1.100 ;
        RECT 267.120 0.820 267.400 1.100 ;
        RECT 268.440 0.820 268.720 1.100 ;
        RECT 270.640 0.820 270.920 1.100 ;
        RECT 271.300 0.820 271.580 1.100 ;
        RECT 271.960 0.820 272.240 1.100 ;
        RECT 272.880 0.820 273.160 1.100 ;
        RECT 273.540 0.820 273.820 1.100 ;
        RECT 274.200 0.820 274.480 1.100 ;
        RECT 275.120 0.820 275.400 1.100 ;
        RECT 275.780 0.820 276.060 1.100 ;
        RECT 276.440 0.820 276.720 1.100 ;
        RECT 277.360 0.820 277.640 1.100 ;
        RECT 278.020 0.820 278.300 1.100 ;
        RECT 278.680 0.820 278.960 1.100 ;
        RECT 279.720 0.820 280.000 1.100 ;
        RECT 280.720 0.820 281.000 1.100 ;
        RECT 281.380 0.820 281.660 1.100 ;
        RECT 282.040 0.820 282.320 1.100 ;
        RECT 282.960 0.820 283.240 1.100 ;
        RECT 283.620 0.820 283.900 1.100 ;
        RECT 284.280 0.820 284.560 1.100 ;
        RECT 285.200 0.820 285.480 1.100 ;
        RECT 285.860 0.820 286.140 1.100 ;
        RECT 286.520 0.820 286.800 1.100 ;
        RECT 287.440 0.820 287.720 1.100 ;
        RECT 288.100 0.820 288.380 1.100 ;
        RECT 288.760 0.820 289.040 1.100 ;
        RECT 289.680 0.820 289.960 1.100 ;
        RECT 290.340 0.820 290.620 1.100 ;
        RECT 291.000 0.820 291.280 1.100 ;
        RECT 291.920 0.820 292.200 1.100 ;
        RECT 292.580 0.820 292.860 1.100 ;
        RECT 293.240 0.820 293.520 1.100 ;
        RECT 294.160 0.820 294.440 1.100 ;
        RECT 294.820 0.820 295.100 1.100 ;
        RECT 295.480 0.820 295.760 1.100 ;
        RECT 296.400 0.820 296.680 1.100 ;
        RECT 297.060 0.820 297.340 1.100 ;
        RECT 297.720 0.820 298.000 1.100 ;
        RECT 298.640 0.820 298.920 1.100 ;
        RECT 299.300 0.820 299.580 1.100 ;
        RECT 299.960 0.820 300.240 1.100 ;
        RECT 301.000 0.820 301.280 1.100 ;
        RECT 302.000 0.820 302.280 1.100 ;
        RECT 302.660 0.820 302.940 1.100 ;
        RECT 303.320 0.820 303.600 1.100 ;
        RECT 304.240 0.820 304.520 1.100 ;
        RECT 304.900 0.820 305.180 1.100 ;
        RECT 305.560 0.820 305.840 1.100 ;
        RECT 306.480 0.820 306.760 1.100 ;
        RECT 307.140 0.820 307.420 1.100 ;
        RECT 307.800 0.820 308.080 1.100 ;
        RECT 308.720 0.820 309.000 1.100 ;
        RECT 309.380 0.820 309.660 1.100 ;
        RECT 310.040 0.820 310.320 1.100 ;
        RECT 310.800 0.820 311.080 1.100 ;
        RECT 312.120 0.820 312.400 1.100 ;
        RECT 314.320 0.820 314.600 1.100 ;
        RECT 314.980 0.820 315.260 1.100 ;
        RECT 315.640 0.820 315.920 1.100 ;
        RECT 316.560 0.820 316.840 1.100 ;
        RECT 317.220 0.820 317.500 1.100 ;
        RECT 317.880 0.820 318.160 1.100 ;
        RECT 318.800 0.820 319.080 1.100 ;
        RECT 319.460 0.820 319.740 1.100 ;
        RECT 320.120 0.820 320.400 1.100 ;
        RECT 321.160 0.820 321.440 1.100 ;
        RECT 322.160 0.820 322.440 1.100 ;
        RECT 322.820 0.820 323.100 1.100 ;
        RECT 323.480 0.820 323.760 1.100 ;
        RECT 324.400 0.820 324.680 1.100 ;
        RECT 325.060 0.820 325.340 1.100 ;
        RECT 325.720 0.820 326.000 1.100 ;
        RECT 326.640 0.820 326.920 1.100 ;
        RECT 327.300 0.820 327.580 1.100 ;
        RECT 327.960 0.820 328.240 1.100 ;
        RECT 328.880 0.820 329.160 1.100 ;
        RECT 329.540 0.820 329.820 1.100 ;
        RECT 330.200 0.820 330.480 1.100 ;
        RECT 331.120 0.820 331.400 1.100 ;
        RECT 331.780 0.820 332.060 1.100 ;
        RECT 332.440 0.820 332.720 1.100 ;
        RECT 333.360 0.820 333.640 1.100 ;
        RECT 334.020 0.820 334.300 1.100 ;
        RECT 334.680 0.820 334.960 1.100 ;
        RECT 335.600 0.820 335.880 1.100 ;
        RECT 336.260 0.820 336.540 1.100 ;
        RECT 336.920 0.820 337.200 1.100 ;
        RECT 337.840 0.820 338.120 1.100 ;
        RECT 338.500 0.820 338.780 1.100 ;
        RECT 339.160 0.820 339.440 1.100 ;
        RECT 340.080 0.820 340.360 1.100 ;
        RECT 340.740 0.820 341.020 1.100 ;
        RECT 341.400 0.820 341.680 1.100 ;
        RECT 342.440 0.820 342.720 1.100 ;
        RECT 343.440 0.820 343.720 1.100 ;
        RECT 344.100 0.820 344.380 1.100 ;
        RECT 344.760 0.820 345.040 1.100 ;
        RECT 345.680 0.820 345.960 1.100 ;
        RECT 346.340 0.820 346.620 1.100 ;
        RECT 347.000 0.820 347.280 1.100 ;
        RECT 347.920 0.820 348.200 1.100 ;
        RECT 348.580 0.820 348.860 1.100 ;
        RECT 349.240 0.820 349.520 1.100 ;
        RECT 350.160 0.820 350.440 1.100 ;
        RECT 350.820 0.820 351.100 1.100 ;
        RECT 351.480 0.820 351.760 1.100 ;
        RECT 352.240 0.820 352.520 1.100 ;
        RECT 353.560 0.820 353.840 1.100 ;
        RECT 355.760 0.820 356.040 1.100 ;
        RECT 356.420 0.820 356.700 1.100 ;
        RECT 357.080 0.820 357.360 1.100 ;
        RECT 358.000 0.820 358.280 1.100 ;
        RECT 358.660 0.820 358.940 1.100 ;
        RECT 359.320 0.820 359.600 1.100 ;
        RECT 360.240 0.820 360.520 1.100 ;
        RECT 360.900 0.820 361.180 1.100 ;
        RECT 361.560 0.820 361.840 1.100 ;
        RECT 362.600 0.820 362.880 1.100 ;
        RECT 363.600 0.820 363.880 1.100 ;
        RECT 364.260 0.820 364.540 1.100 ;
        RECT 364.920 0.820 365.200 1.100 ;
        RECT 365.840 0.820 366.120 1.100 ;
        RECT 366.500 0.820 366.780 1.100 ;
        RECT 367.160 0.820 367.440 1.100 ;
        RECT 368.080 0.820 368.360 1.100 ;
        RECT 368.740 0.820 369.020 1.100 ;
        RECT 369.400 0.820 369.680 1.100 ;
        RECT 370.320 0.820 370.600 1.100 ;
        RECT 370.980 0.820 371.260 1.100 ;
        RECT 371.640 0.820 371.920 1.100 ;
        RECT 372.560 0.820 372.840 1.100 ;
        RECT 373.220 0.820 373.500 1.100 ;
        RECT 373.880 0.820 374.160 1.100 ;
        RECT 374.800 0.820 375.080 1.100 ;
        RECT 375.460 0.820 375.740 1.100 ;
        RECT 376.120 0.820 376.400 1.100 ;
        RECT 377.040 0.820 377.320 1.100 ;
        RECT 377.700 0.820 377.980 1.100 ;
        RECT 378.360 0.820 378.640 1.100 ;
        RECT 379.280 0.820 379.560 1.100 ;
        RECT 379.940 0.820 380.220 1.100 ;
        RECT 380.600 0.820 380.880 1.100 ;
        RECT 381.520 0.820 381.800 1.100 ;
        RECT 382.180 0.820 382.460 1.100 ;
        RECT 382.840 0.820 383.120 1.100 ;
        RECT 383.880 0.820 384.160 1.100 ;
        RECT 384.880 0.820 385.160 1.100 ;
        RECT 385.540 0.820 385.820 1.100 ;
        RECT 386.200 0.820 386.480 1.100 ;
        RECT 387.120 0.820 387.400 1.100 ;
        RECT 387.780 0.820 388.060 1.100 ;
        RECT 388.440 0.820 388.720 1.100 ;
        RECT 389.360 0.820 389.640 1.100 ;
        RECT 390.020 0.820 390.300 1.100 ;
        RECT 390.680 0.820 390.960 1.100 ;
        RECT 391.600 0.820 391.880 1.100 ;
        RECT 392.260 0.820 392.540 1.100 ;
        RECT 392.920 0.820 393.200 1.100 ;
        RECT 393.840 0.820 394.120 1.100 ;
        RECT 394.500 0.820 394.780 1.100 ;
        RECT 395.160 0.820 395.440 1.100 ;
        RECT 395.920 0.820 396.200 1.100 ;
        RECT 397.240 0.820 397.520 1.100 ;
        RECT 399.440 0.820 399.720 1.100 ;
        RECT 400.100 0.820 400.380 1.100 ;
        RECT 400.760 0.820 401.040 1.100 ;
        RECT 401.680 0.820 401.960 1.100 ;
        RECT 402.340 0.820 402.620 1.100 ;
        RECT 403.000 0.820 403.280 1.100 ;
        RECT 404.040 0.820 404.320 1.100 ;
        RECT 405.040 0.820 405.320 1.100 ;
        RECT 405.700 0.820 405.980 1.100 ;
        RECT 406.360 0.820 406.640 1.100 ;
        RECT 407.280 0.820 407.560 1.100 ;
        RECT 407.940 0.820 408.220 1.100 ;
        RECT 408.600 0.820 408.880 1.100 ;
        RECT 409.520 0.820 409.800 1.100 ;
        RECT 410.180 0.820 410.460 1.100 ;
        RECT 410.840 0.820 411.120 1.100 ;
        RECT 411.760 0.820 412.040 1.100 ;
        RECT 412.420 0.820 412.700 1.100 ;
        RECT 413.080 0.820 413.360 1.100 ;
        RECT 414.000 0.820 414.280 1.100 ;
        RECT 414.660 0.820 414.940 1.100 ;
        RECT 415.320 0.820 415.600 1.100 ;
        RECT 416.240 0.820 416.520 1.100 ;
        RECT 416.900 0.820 417.180 1.100 ;
        RECT 417.560 0.820 417.840 1.100 ;
        RECT 418.480 0.820 418.760 1.100 ;
        RECT 419.140 0.820 419.420 1.100 ;
        RECT 419.800 0.820 420.080 1.100 ;
        RECT 420.720 0.820 421.000 1.100 ;
        RECT 421.380 0.820 421.660 1.100 ;
        RECT 422.040 0.820 422.320 1.100 ;
        RECT 422.960 0.820 423.240 1.100 ;
        RECT 423.620 0.820 423.900 1.100 ;
        RECT 424.280 0.820 424.560 1.100 ;
        RECT 425.320 0.820 425.600 1.100 ;
        RECT 426.320 0.820 426.600 1.100 ;
        RECT 426.980 0.820 427.260 1.100 ;
        RECT 427.640 0.820 427.920 1.100 ;
        RECT 428.560 0.820 428.840 1.100 ;
        RECT 429.220 0.820 429.500 1.100 ;
        RECT 429.880 0.820 430.160 1.100 ;
        RECT 430.800 0.820 431.080 1.100 ;
        RECT 431.460 0.820 431.740 1.100 ;
        RECT 432.120 0.820 432.400 1.100 ;
        RECT 433.040 0.820 433.320 1.100 ;
        RECT 433.700 0.820 433.980 1.100 ;
        RECT 434.360 0.820 434.640 1.100 ;
        RECT 435.280 0.820 435.560 1.100 ;
        RECT 435.940 0.820 436.220 1.100 ;
        RECT 436.600 0.820 436.880 1.100 ;
        RECT 437.360 0.820 437.640 1.100 ;
        RECT 438.680 0.820 438.960 1.100 ;
        RECT 440.880 0.820 441.160 1.100 ;
        RECT 441.540 0.820 441.820 1.100 ;
        RECT 442.200 0.820 442.480 1.100 ;
        RECT 443.120 0.820 443.400 1.100 ;
        RECT 443.780 0.820 444.060 1.100 ;
        RECT 444.440 0.820 444.720 1.100 ;
        RECT 445.480 0.820 445.760 1.100 ;
        RECT 446.480 0.820 446.760 1.100 ;
        RECT 447.140 0.820 447.420 1.100 ;
        RECT 447.800 0.820 448.080 1.100 ;
        RECT 448.720 0.820 449.000 1.100 ;
        RECT 449.380 0.820 449.660 1.100 ;
        RECT 450.040 0.820 450.320 1.100 ;
        RECT 450.960 0.820 451.240 1.100 ;
        RECT 451.620 0.820 451.900 1.100 ;
        RECT 452.280 0.820 452.560 1.100 ;
        RECT 453.200 0.820 453.480 1.100 ;
        RECT 453.860 0.820 454.140 1.100 ;
        RECT 454.520 0.820 454.800 1.100 ;
        RECT 455.440 0.820 455.720 1.100 ;
        RECT 456.100 0.820 456.380 1.100 ;
        RECT 456.760 0.820 457.040 1.100 ;
        RECT 457.680 0.820 457.960 1.100 ;
        RECT 458.340 0.820 458.620 1.100 ;
        RECT 459.000 0.820 459.280 1.100 ;
        RECT 459.920 0.820 460.200 1.100 ;
        RECT 460.580 0.820 460.860 1.100 ;
        RECT 461.240 0.820 461.520 1.100 ;
        RECT 462.160 0.820 462.440 1.100 ;
        RECT 462.820 0.820 463.100 1.100 ;
        RECT 463.480 0.820 463.760 1.100 ;
        RECT 464.400 0.820 464.680 1.100 ;
        RECT 465.060 0.820 465.340 1.100 ;
        RECT 465.720 0.820 466.000 1.100 ;
        RECT 466.760 0.820 467.040 1.100 ;
        RECT 467.760 0.820 468.040 1.100 ;
        RECT 468.420 0.820 468.700 1.100 ;
        RECT 469.080 0.820 469.360 1.100 ;
        RECT 470.000 0.820 470.280 1.100 ;
        RECT 470.660 0.820 470.940 1.100 ;
        RECT 471.320 0.820 471.600 1.100 ;
        RECT 472.240 0.820 472.520 1.100 ;
        RECT 472.900 0.820 473.180 1.100 ;
        RECT 473.560 0.820 473.840 1.100 ;
        RECT 474.480 0.820 474.760 1.100 ;
        RECT 475.140 0.820 475.420 1.100 ;
        RECT 475.800 0.820 476.080 1.100 ;
        RECT 476.720 0.820 477.000 1.100 ;
        RECT 477.380 0.820 477.660 1.100 ;
        RECT 478.040 0.820 478.320 1.100 ;
        RECT 478.960 0.820 479.240 1.100 ;
        RECT 479.620 0.820 479.900 1.100 ;
        RECT 480.280 0.820 480.560 1.100 ;
        RECT 481.040 0.820 481.320 1.100 ;
        RECT 482.360 0.820 482.640 1.100 ;
        RECT 484.560 0.820 484.840 1.100 ;
        RECT 485.220 0.820 485.500 1.100 ;
        RECT 485.880 0.820 486.160 1.100 ;
        RECT 486.920 0.820 487.200 1.100 ;
        RECT 487.920 0.820 488.200 1.100 ;
        RECT 488.580 0.820 488.860 1.100 ;
        RECT 489.240 0.820 489.520 1.100 ;
        RECT 490.160 0.820 490.440 1.100 ;
        RECT 490.820 0.820 491.100 1.100 ;
        RECT 491.480 0.820 491.760 1.100 ;
        RECT 492.400 0.820 492.680 1.100 ;
        RECT 493.060 0.820 493.340 1.100 ;
        RECT 493.720 0.820 494.000 1.100 ;
        RECT 494.640 0.820 494.920 1.100 ;
        RECT 495.300 0.820 495.580 1.100 ;
        RECT 495.960 0.820 496.240 1.100 ;
        RECT 496.880 0.820 497.160 1.100 ;
        RECT 497.540 0.820 497.820 1.100 ;
        RECT 498.200 0.820 498.480 1.100 ;
        RECT 499.120 0.820 499.400 1.100 ;
        RECT 499.780 0.820 500.060 1.100 ;
        RECT 500.440 0.820 500.720 1.100 ;
        RECT 501.360 0.820 501.640 1.100 ;
        RECT 502.020 0.820 502.300 1.100 ;
        RECT 502.680 0.820 502.960 1.100 ;
        RECT 503.600 0.820 503.880 1.100 ;
        RECT 504.260 0.820 504.540 1.100 ;
        RECT 504.920 0.820 505.200 1.100 ;
        RECT 505.840 0.820 506.120 1.100 ;
        RECT 506.500 0.820 506.780 1.100 ;
        RECT 507.160 0.820 507.440 1.100 ;
        RECT 508.200 0.820 508.480 1.100 ;
        RECT 509.200 0.820 509.480 1.100 ;
        RECT 509.860 0.820 510.140 1.100 ;
        RECT 510.520 0.820 510.800 1.100 ;
        RECT 511.440 0.820 511.720 1.100 ;
        RECT 512.100 0.820 512.380 1.100 ;
        RECT 512.760 0.820 513.040 1.100 ;
        RECT 513.680 0.820 513.960 1.100 ;
        RECT 514.340 0.820 514.620 1.100 ;
        RECT 515.000 0.820 515.280 1.100 ;
        RECT 515.920 0.820 516.200 1.100 ;
        RECT 516.580 0.820 516.860 1.100 ;
        RECT 517.240 0.820 517.520 1.100 ;
        RECT 518.160 0.820 518.440 1.100 ;
        RECT 518.820 0.820 519.100 1.100 ;
        RECT 519.480 0.820 519.760 1.100 ;
        RECT 520.400 0.820 520.680 1.100 ;
        RECT 521.060 0.820 521.340 1.100 ;
        RECT 521.720 0.820 522.000 1.100 ;
        RECT 522.480 0.820 522.760 1.100 ;
        RECT 523.800 0.820 524.080 1.100 ;
        RECT 526.000 0.820 526.280 1.100 ;
        RECT 526.660 0.820 526.940 1.100 ;
        RECT 527.320 0.820 527.600 1.100 ;
        RECT 528.360 0.820 528.640 1.100 ;
        RECT 529.360 0.820 529.640 1.100 ;
        RECT 530.020 0.820 530.300 1.100 ;
        RECT 530.680 0.820 530.960 1.100 ;
        RECT 531.600 0.820 531.880 1.100 ;
        RECT 532.260 0.820 532.540 1.100 ;
        RECT 532.920 0.820 533.200 1.100 ;
        RECT 533.840 0.820 534.120 1.100 ;
        RECT 534.500 0.820 534.780 1.100 ;
        RECT 535.160 0.820 535.440 1.100 ;
        RECT 536.080 0.820 536.360 1.100 ;
        RECT 536.740 0.820 537.020 1.100 ;
        RECT 537.400 0.820 537.680 1.100 ;
        RECT 538.320 0.820 538.600 1.100 ;
        RECT 538.980 0.820 539.260 1.100 ;
        RECT 539.640 0.820 539.920 1.100 ;
        RECT 540.560 0.820 540.840 1.100 ;
        RECT 541.220 0.820 541.500 1.100 ;
        RECT 541.880 0.820 542.160 1.100 ;
        RECT 542.800 0.820 543.080 1.100 ;
        RECT 543.460 0.820 543.740 1.100 ;
        RECT 544.120 0.820 544.400 1.100 ;
        RECT 545.040 0.820 545.320 1.100 ;
        RECT 545.700 0.820 545.980 1.100 ;
        RECT 546.360 0.820 546.640 1.100 ;
        RECT 547.280 0.820 547.560 1.100 ;
        RECT 547.940 0.820 548.220 1.100 ;
        RECT 548.600 0.820 548.880 1.100 ;
        RECT 549.640 0.820 549.920 1.100 ;
        RECT 550.640 0.820 550.920 1.100 ;
        RECT 551.300 0.820 551.580 1.100 ;
        RECT 551.960 0.820 552.240 1.100 ;
        RECT 552.880 0.820 553.160 1.100 ;
        RECT 553.540 0.820 553.820 1.100 ;
        RECT 554.200 0.820 554.480 1.100 ;
        RECT 555.120 0.820 555.400 1.100 ;
        RECT 555.780 0.820 556.060 1.100 ;
        RECT 556.440 0.820 556.720 1.100 ;
        RECT 557.360 0.820 557.640 1.100 ;
        RECT 558.020 0.820 558.300 1.100 ;
        RECT 558.680 0.820 558.960 1.100 ;
        RECT 559.600 0.820 559.880 1.100 ;
        RECT 560.260 0.820 560.540 1.100 ;
        RECT 560.920 0.820 561.200 1.100 ;
        RECT 561.840 0.820 562.120 1.100 ;
        RECT 562.500 0.820 562.780 1.100 ;
        RECT 563.160 0.820 563.440 1.100 ;
        RECT 564.080 0.820 564.360 1.100 ;
        RECT 564.740 0.820 565.020 1.100 ;
        RECT 565.400 0.820 565.680 1.100 ;
        RECT 566.160 0.820 566.440 1.100 ;
        RECT 567.480 0.820 567.760 1.100 ;
        RECT 569.800 0.820 570.080 1.100 ;
        RECT 570.800 0.820 571.080 1.100 ;
        RECT 571.460 0.820 571.740 1.100 ;
        RECT 572.120 0.820 572.400 1.100 ;
        RECT 573.040 0.820 573.320 1.100 ;
        RECT 573.700 0.820 573.980 1.100 ;
        RECT 574.360 0.820 574.640 1.100 ;
        RECT 575.280 0.820 575.560 1.100 ;
        RECT 575.940 0.820 576.220 1.100 ;
        RECT 576.600 0.820 576.880 1.100 ;
        RECT 577.520 0.820 577.800 1.100 ;
        RECT 578.180 0.820 578.460 1.100 ;
        RECT 578.840 0.820 579.120 1.100 ;
        RECT 579.760 0.820 580.040 1.100 ;
        RECT 580.420 0.820 580.700 1.100 ;
        RECT 581.080 0.820 581.360 1.100 ;
        RECT 582.000 0.820 582.280 1.100 ;
        RECT 582.660 0.820 582.940 1.100 ;
        RECT 583.320 0.820 583.600 1.100 ;
        RECT 584.240 0.820 584.520 1.100 ;
        RECT 584.900 0.820 585.180 1.100 ;
        RECT 585.560 0.820 585.840 1.100 ;
        RECT 586.480 0.820 586.760 1.100 ;
        RECT 587.140 0.820 587.420 1.100 ;
        RECT 587.800 0.820 588.080 1.100 ;
        RECT 588.720 0.820 589.000 1.100 ;
        RECT 589.380 0.820 589.660 1.100 ;
        RECT 590.040 0.820 590.320 1.100 ;
        RECT 591.080 0.820 591.360 1.100 ;
        RECT 592.080 0.820 592.360 1.100 ;
        RECT 592.740 0.820 593.020 1.100 ;
        RECT 593.400 0.820 593.680 1.100 ;
        RECT 594.320 0.820 594.600 1.100 ;
        RECT 594.980 0.820 595.260 1.100 ;
        RECT 595.640 0.820 595.920 1.100 ;
        RECT 596.560 0.820 596.840 1.100 ;
        RECT 597.220 0.820 597.500 1.100 ;
        RECT 597.880 0.820 598.160 1.100 ;
        RECT 598.800 0.820 599.080 1.100 ;
        RECT 599.460 0.820 599.740 1.100 ;
        RECT 600.120 0.820 600.400 1.100 ;
        RECT 601.040 0.820 601.320 1.100 ;
        RECT 601.700 0.820 601.980 1.100 ;
        RECT 602.360 0.820 602.640 1.100 ;
        RECT 603.280 0.820 603.560 1.100 ;
        RECT 603.940 0.820 604.220 1.100 ;
        RECT 604.600 0.820 604.880 1.100 ;
        RECT 605.520 0.820 605.800 1.100 ;
        RECT 606.180 0.820 606.460 1.100 ;
        RECT 606.840 0.820 607.120 1.100 ;
        RECT 607.600 0.820 607.880 1.100 ;
        RECT 608.920 0.820 609.200 1.100 ;
        RECT 611.240 0.820 611.520 1.100 ;
        RECT 612.240 0.820 612.520 1.100 ;
        RECT 612.900 0.820 613.180 1.100 ;
        RECT 613.560 0.820 613.840 1.100 ;
        RECT 614.480 0.820 614.760 1.100 ;
        RECT 615.140 0.820 615.420 1.100 ;
        RECT 615.800 0.820 616.080 1.100 ;
        RECT 616.720 0.820 617.000 1.100 ;
        RECT 617.380 0.820 617.660 1.100 ;
        RECT 618.040 0.820 618.320 1.100 ;
        RECT 618.960 0.820 619.240 1.100 ;
        RECT 619.620 0.820 619.900 1.100 ;
        RECT 620.280 0.820 620.560 1.100 ;
        RECT 621.200 0.820 621.480 1.100 ;
        RECT 621.860 0.820 622.140 1.100 ;
        RECT 622.520 0.820 622.800 1.100 ;
        RECT 623.440 0.820 623.720 1.100 ;
        RECT 624.100 0.820 624.380 1.100 ;
        RECT 624.760 0.820 625.040 1.100 ;
        RECT 625.680 0.820 625.960 1.100 ;
        RECT 626.340 0.820 626.620 1.100 ;
        RECT 627.000 0.820 627.280 1.100 ;
        RECT 627.920 0.820 628.200 1.100 ;
        RECT 628.580 0.820 628.860 1.100 ;
        RECT 629.240 0.820 629.520 1.100 ;
        RECT 630.160 0.820 630.440 1.100 ;
        RECT 630.820 0.820 631.100 1.100 ;
        RECT 631.480 0.820 631.760 1.100 ;
        RECT 632.520 0.820 632.800 1.100 ;
        RECT 633.520 0.820 633.800 1.100 ;
        RECT 634.180 0.820 634.460 1.100 ;
        RECT 634.840 0.820 635.120 1.100 ;
        RECT 635.760 0.820 636.040 1.100 ;
        RECT 636.420 0.820 636.700 1.100 ;
        RECT 637.080 0.820 637.360 1.100 ;
        RECT 638.000 0.820 638.280 1.100 ;
        RECT 638.660 0.820 638.940 1.100 ;
        RECT 639.320 0.820 639.600 1.100 ;
        RECT 640.240 0.820 640.520 1.100 ;
        RECT 640.900 0.820 641.180 1.100 ;
        RECT 641.560 0.820 641.840 1.100 ;
        RECT 642.480 0.820 642.760 1.100 ;
        RECT 643.140 0.820 643.420 1.100 ;
        RECT 643.800 0.820 644.080 1.100 ;
        RECT 644.720 0.820 645.000 1.100 ;
        RECT 645.380 0.820 645.660 1.100 ;
        RECT 646.040 0.820 646.320 1.100 ;
        RECT 646.960 0.820 647.240 1.100 ;
        RECT 647.620 0.820 647.900 1.100 ;
        RECT 648.280 0.820 648.560 1.100 ;
        RECT 649.200 0.820 649.480 1.100 ;
        RECT 649.860 0.820 650.140 1.100 ;
        RECT 650.520 0.820 650.800 1.100 ;
        RECT 651.280 0.820 651.560 1.100 ;
        RECT 652.600 0.820 652.880 1.100 ;
        RECT 654.920 0.820 655.200 1.100 ;
        RECT 655.920 0.820 656.200 1.100 ;
        RECT 656.580 0.820 656.860 1.100 ;
        RECT 657.240 0.820 657.520 1.100 ;
        RECT 658.160 0.820 658.440 1.100 ;
        RECT 658.820 0.820 659.100 1.100 ;
        RECT 659.480 0.820 659.760 1.100 ;
        RECT 660.400 0.820 660.680 1.100 ;
        RECT 661.060 0.820 661.340 1.100 ;
        RECT 661.720 0.820 662.000 1.100 ;
        RECT 662.640 0.820 662.920 1.100 ;
        RECT 663.300 0.820 663.580 1.100 ;
        RECT 663.960 0.820 664.240 1.100 ;
        RECT 664.880 0.820 665.160 1.100 ;
        RECT 665.540 0.820 665.820 1.100 ;
        RECT 666.200 0.820 666.480 1.100 ;
        RECT 667.120 0.820 667.400 1.100 ;
        RECT 667.780 0.820 668.060 1.100 ;
        RECT 668.440 0.820 668.720 1.100 ;
        RECT 669.360 0.820 669.640 1.100 ;
        RECT 670.020 0.820 670.300 1.100 ;
        RECT 670.680 0.820 670.960 1.100 ;
        RECT 671.600 0.820 671.880 1.100 ;
        RECT 672.260 0.820 672.540 1.100 ;
        RECT 672.920 0.820 673.200 1.100 ;
        RECT 673.840 0.820 674.120 1.100 ;
        RECT 674.500 0.820 674.780 1.100 ;
        RECT 675.160 0.820 675.440 1.100 ;
        RECT 676.200 0.820 676.480 1.100 ;
        RECT 677.200 0.820 677.480 1.100 ;
        RECT 677.860 0.820 678.140 1.100 ;
        RECT 678.520 0.820 678.800 1.100 ;
        RECT 679.540 0.820 679.820 1.100 ;
      LAYER Metal4 ;
        RECT 4.610 47.805 4.990 48.185 ;
        RECT 4.635 47.525 4.965 47.805 ;
        RECT 4.610 47.145 4.990 47.525 ;
        RECT 4.635 46.865 4.965 47.145 ;
        RECT 4.610 46.485 4.990 46.865 ;
        RECT 4.635 8.470 4.965 46.485 ;
        RECT 53.580 45.105 53.960 45.485 ;
        RECT 53.605 44.825 53.935 45.105 ;
        RECT 53.580 44.445 53.960 44.825 ;
        RECT 53.605 44.165 53.935 44.445 ;
        RECT 53.580 43.785 53.960 44.165 ;
        RECT 38.750 24.905 39.130 25.285 ;
        RECT 38.775 24.625 39.105 24.905 ;
        RECT 38.750 24.245 39.130 24.625 ;
        RECT 38.775 23.965 39.105 24.245 ;
        RECT 38.750 23.585 39.130 23.965 ;
        RECT 22.800 22.205 23.180 22.585 ;
        RECT 22.825 21.925 23.155 22.205 ;
        RECT 22.800 21.545 23.180 21.925 ;
        RECT 22.825 21.265 23.155 21.545 ;
        RECT 22.800 20.885 23.180 21.265 ;
        RECT 22.825 8.470 23.155 20.885 ;
        RECT 38.775 8.470 39.105 23.585 ;
        RECT 53.605 8.470 53.935 43.785 ;
        RECT 72.890 42.405 73.270 42.785 ;
        RECT 72.915 42.125 73.245 42.405 ;
        RECT 72.890 41.745 73.270 42.125 ;
        RECT 72.915 41.465 73.245 41.745 ;
        RECT 72.890 41.085 73.270 41.465 ;
        RECT 72.915 8.470 73.245 41.085 ;
        RECT 121.860 39.705 122.240 40.085 ;
        RECT 121.885 39.425 122.215 39.705 ;
        RECT 121.860 39.045 122.240 39.425 ;
        RECT 121.885 38.765 122.215 39.045 ;
        RECT 121.860 38.385 122.240 38.765 ;
        RECT 107.030 30.305 107.410 30.685 ;
        RECT 107.055 30.025 107.385 30.305 ;
        RECT 107.030 29.645 107.410 30.025 ;
        RECT 107.055 29.365 107.385 29.645 ;
        RECT 107.030 28.985 107.410 29.365 ;
        RECT 87.720 27.605 88.100 27.985 ;
        RECT 87.745 27.325 88.075 27.605 ;
        RECT 87.720 26.945 88.100 27.325 ;
        RECT 87.745 26.665 88.075 26.945 ;
        RECT 87.720 26.285 88.100 26.665 ;
        RECT 87.745 8.470 88.075 26.285 ;
        RECT 107.055 8.470 107.385 28.985 ;
        RECT 121.885 8.470 122.215 38.385 ;
        RECT 4.610 8.090 4.990 8.470 ;
        RECT 22.800 8.090 23.180 8.470 ;
        RECT 38.750 8.090 39.130 8.470 ;
        RECT 53.580 8.090 53.960 8.470 ;
        RECT 72.890 8.090 73.270 8.470 ;
        RECT 87.720 8.090 88.100 8.470 ;
        RECT 107.030 8.090 107.410 8.470 ;
        RECT 121.860 8.090 122.240 8.470 ;
        RECT 4.635 7.810 4.965 8.090 ;
        RECT 22.825 7.810 23.155 8.090 ;
        RECT 38.775 7.810 39.105 8.090 ;
        RECT 53.605 7.810 53.935 8.090 ;
        RECT 72.915 7.810 73.245 8.090 ;
        RECT 87.745 7.810 88.075 8.090 ;
        RECT 107.055 7.810 107.385 8.090 ;
        RECT 121.885 7.810 122.215 8.090 ;
        RECT 4.610 7.430 4.990 7.810 ;
        RECT 22.800 7.430 23.180 7.810 ;
        RECT 38.750 7.430 39.130 7.810 ;
        RECT 53.580 7.430 53.960 7.810 ;
        RECT 72.890 7.430 73.270 7.810 ;
        RECT 87.720 7.430 88.100 7.810 ;
        RECT 107.030 7.430 107.410 7.810 ;
        RECT 121.860 7.430 122.240 7.810 ;
        RECT 4.635 7.150 4.965 7.430 ;
        RECT 22.825 7.150 23.155 7.430 ;
        RECT 38.775 7.150 39.105 7.430 ;
        RECT 53.605 7.150 53.935 7.430 ;
        RECT 72.915 7.150 73.245 7.430 ;
        RECT 87.745 7.150 88.075 7.430 ;
        RECT 107.055 7.150 107.385 7.430 ;
        RECT 121.885 7.150 122.215 7.430 ;
        RECT 4.610 6.770 4.990 7.150 ;
        RECT 22.800 6.770 23.180 7.150 ;
        RECT 38.750 6.770 39.130 7.150 ;
        RECT 53.580 6.770 53.960 7.150 ;
        RECT 72.890 6.770 73.270 7.150 ;
        RECT 87.720 6.770 88.100 7.150 ;
        RECT 107.030 6.770 107.410 7.150 ;
        RECT 121.860 6.770 122.240 7.150 ;
  END
END efuse_array
END LIBRARY

