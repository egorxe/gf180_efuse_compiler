.option TEMP=25.0

.include "design.xyce"
.lib "sm141064.xyce" typical
.lib "sm141064.xyce" efuse
.lib "sm141064.xyce" diode_typical

.include efuse_ctrl.spice

Xtest wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[1] wb_adr_i[2]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[1] wb_dat_i[2] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5]
+ wb_dat_i[6] wb_dat_i[7] wb_dat_o[0] wb_dat_o[1] wb_dat_o[2] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_rst_i wb_sel_i wb_stb_i wb_we_i VDD VSS efuse_ctrl


VGND GND 0 0V
VVDD VDD GND 5V ;PULSE(0 5V 2ns 1ns 1ns 8ms 20ms)
VVSS VSS GND 0V

* WB test
Vadr[0] wb_adr_i[0] 0 PWL 0ns 0V 50ns 0V 51ns 5V
Vadr[1] wb_adr_i[1] 0 0V
Vadr[2] wb_adr_i[2] 0 5V
Vadr[3] wb_adr_i[3] 0 0V
Vadr[4] wb_adr_i[4] 0 0V
Vadr[5] wb_adr_i[5] 0 0V
Vadr[6] wb_adr_i[6] 0 5V
Vadr[7] wb_adr_i[7] 0 5V
Vadr[8] wb_adr_i[8] 0 5V
Vadr[9] wb_adr_i[9] 0 0V
Vadr[10] wb_adr_i[10] 0 0V
Vadr[11] wb_adr_i[11] 0 PWL 0ns 0V 30.9ns 0V 31ns 5V 50.9ns 5V 51ns 0V

Vdat[0] wb_dat_i[0] 0 5V
Vdat[1] wb_dat_i[1] 0 0V
Vdat[2] wb_dat_i[2] 0 0V
Vdat[3] wb_dat_i[3] 0 0V
Vdat[4] wb_dat_i[4] 0 5V
Vdat[5] wb_dat_i[5] 0 0V
Vdat[6] wb_dat_i[6] 0 0V
Vdat[7] wb_dat_i[7] 0 0V

Vclk wb_clk_i GND PULSE(0 5V 0us 0.1ns 0.1ns 10ns 20ns)

Vwe wb_we_i GND 0 PWL 0ns 0V 30.9ns 0V 31ns 5V 50.9ns 5V 51ns 0V

Vrst wb_rst_i GND PWL 0ns 5V 10.9ns 5V 11ns 0V
Vstb wb_stb_i GND PWL 0ns 0V 30.9ns 0V 31ns 5V 50.9ns 5V 51ns 0V 70.9ns 0V 71ns 5V 90.9ns 5V 91ns 0V


.TRAN 1e-9 300e-9 UIC
.PRINT TRAN V(wb_clk_i) V(wb_rst_i) V(wb_stb_i) V(wb_dat_o[0]) V(wb_dat_o[1]) V(wb_dat_o[2]) V(wb_dat_o[3]) V(wb_dat_o[4]) V(wb_dat_o[5]) V(wb_dat_o[6]) V(wb_dat_o[7]) V(wb_ack_o) 
+ I(XTEST:Xefuse_array*:X*:RFUSE*)

.end

