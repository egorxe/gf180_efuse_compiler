.option TEMP=25.0

.include "design.xyce"
.lib "sm141064.xyce" typical
.lib "sm141064.xyce" efuse

.include efuse_array.spice

Xtest COL_PROG[0] COL_PROG[1] COL_PROG[2] COL_PROG[3] COL_PROG[4] COL_PROG[5]
+ COL_PROG[6] COL_PROG[7] DO[0] LINE[0] DO[1] DO[2] DO[3] LINE[1] DO[4] DO[5] LINE[2]
+ DO[6] DO[7] LINE[3] LINE[4] LINE[5] LINE[6] LINE[7] LINE[8] LINE[9] LINE[10] LINE[11]
+ LINE[12] LINE[13] LINE[14] LINE[15] SENSE nPRESET VSS VDD efuse_array


VGND GND 0 0V
VVDD VDD GND 5V
VVSS VSS GND 0V

* programming test
VLINE[0] LINE[0] GND 0
VLINE[1] LINE[1] GND 0
VLINE[2] LINE[2] GND 0V
VLINE[3] LINE[3] GND 5V
VLINE[4] LINE[4] GND 0
VLINE[5] LINE[5] GND 0
VLINE[6] LINE[6] GND 0
VLINE[7] LINE[7] GND 0
VLINE[8] LINE[8] GND 0
VLINE[9] LINE[9] GND 0
VLINE[10] LINE[10] GND 0
VLINE[11] LINE[11] GND 0
VLINE[12] LINE[12] GND 0
VLINE[13] LINE[13] GND 0
VLINE[14] LINE[14] GND 0
VLINE[15] LINE[15] GND 0

*VCOL1_PROG COL_PROG[1] GND 5V
VCOL2_PROG COL_PROG[2] GND 5V
VCOL3_PROG COL_PROG[3] GND 5V
VCOL4_PROG COL_PROG[4] GND 5V
VCOL5_PROG COL_PROG[5] GND 5V
VCOL6_PROG COL_PROG[6] GND 5V
VCOL7_PROG COL_PROG[7] GND 5V

VCOL0_PROG COL_PROG[0] GND PULSE(5V 0V 1us 10ns 10ns 100ns 100us)
VCOL1_PROG COL_PROG[1] GND PULSE(5V 0V 1us 10ns 10ns 100ns 100us)
VPRESET nPRESET GND 5V
VSENSE SENSE GND 0

* sense test
*VCOL0_PROG COL_PROG[0] GND 5V
*VPRESET nPRESET GND PULSE(5V 0V 1020ns 1ns 1ns 10ns 100us)
*VSENSE SENSE GND PULSE(0 5V 1050ns 1ns 1ns 10ns 10us)



.TRAN 1e-12 1.5e-6
.PRINT TRAN V(DO[0]) V(DO[1]) V(DO[2]) V(DO[3]) V(DO[4]) V(DO[5]) V(DO[6]) V(DO[7]) V(nPRESET) V(COL_PROG[0])
+I(VVDD) I(XTEST:X*:RFUSE*)
.end

